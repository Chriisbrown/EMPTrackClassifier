library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_misc.all;
  use ieee.numeric_std.all;

  use work.Constants.all;
  use work.Types.all;
  package Arrays0 is

    constant initPredict : ty := to_ty(0);
    constant feature : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((4, 1, 0, 0, 1, 0, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 1, 0, 0, 19, 2, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 1, 0, 3, 1, 2, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 4, 4, 4, 3, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 4, 4, 4, 16, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 4, 4, 3, 17, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 1, 0, 0, 19, 2, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 4, 4, 4, 1, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 3, 0, 17, 1, 2, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 4, 4, 4, 17, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 1, 4, 3, 0, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 16, 0, 1, 3, 2, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 4, 4, 17, 2, 17, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 1, 4, 4, 0, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 2, 4, 1, 17, 17, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 2, 4, 3, 17, 17, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 4, 1, 10, 2, 3, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 16, 2, 10, 18, 3, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 1, 4, 18, 4, 20, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 1, 4, 18, 3, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 2, 1, 4, 17, 3, 12, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 2, 1, 3, 0, 18, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 18, 2, 4, 18, 16, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 4, 4, 10, 2, 20, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 2, 1, 18, 7, 4, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 1, 2, 18, 17, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 4, 1, 0, 2, 18, 12, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 18, 1, 18, 4, 5, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 18, 4, 1, 4, 17, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 18, 1, 18, 4, 16, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 2, 16, 3, 7, 17, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 17, 2, 5, 16, 3, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (7, 17, 6, 5, 12, 20, 13, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 7, 18, 17, 6, 4, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 7, 3, 17, 6, 14, 14, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 4, 18, 0, 16, 4, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 1, 16, 17, 16, -2, 12, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 7, 16, 13, 6, 20, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 18, 18, -2, 18, 18, 20, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 2, 17, 7, 18, 7, 12, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 5, 17, 8, 2, 7, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 17, 2, 7, 13, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 20, 16, 10, 16, 20, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 4, 18, 19, 1, 3, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 1, 17, 5, 16, -2, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 17, 17, 4, 17, 7, 12, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 5, 18, 8, 2, 4, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 3, 3, 18, 2, 16, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 20, 17, 17, 16, 7, 12, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 1, 16, 0, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 17, 8, 7, 15, 13, 5, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 5, 17, 8, 14, 7, 12, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 3, 16, 18, 2, -2, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 18, 4, 18, 3, 19, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 6, 1, -2, 7, 2, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 18, 20, 18, 5, 19, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 1, 4, 5, 17, 1, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 20, 16, 10, 16, 16, 10, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 6, 18, -2, 7, 3, 20, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 2, 17, 6, 17, 7, 12, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 20, 4, 10, 2, 1, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 5, 16, 8, 17, 1, 19, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 17, 8, 7, 12, 13, 5, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 19, 3, 6, 17, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 3, 4, 18, 2, 2, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 18, 20, 4, 4, 19, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 1, 16, 0, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 19, 16, 6, 17, 2, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 6, 19, 4, 2, 11, 12, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 5, 17, 17, 16, 6, 14, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 18, 16, 18, 20, 17, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, -2, 3, 17, 3, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 5, 19, 7, 4, 10, 12, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 2, 17, 4, -2, 7, 14, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 7, 14, 5, 13, 15, 13, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 4, 17, 16, 16, 7, 14, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 18, 4, 4, 1, 2, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 18, -2, 3, 3, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 0, 17, 18, 3, -2, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 4, 0, 5, 16, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 0, 4, 2, 5, 17, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 19, 3, 20, -2, 2, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 3, 4, 4, 19, 18, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 13, 13, 7, 19, 15, 12, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 6, 17, 4, 3, 2, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (15, 17, 17, 13, 14, 12, 13, -2, -2, -2, -2, -2, -2, -2, -2),
                (5, 8, 17, 17, 7, 4, 10, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 3, -2, 1, 3, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 16, 4, 2, 15, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 8, 17, 2, 5, 2, 10, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 15, -2, 20, 17, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 18, 4, 4, 4, 20, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 3, 16, 4, 1, -2, 14, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 3, 4, 1, 1, 1, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 2, -2, 7, 10, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 20, 11, -2, -2, 2, 19, -2, -2, -2, -2, -2, -2, -2, -2),
                (5, 16, 2, 2, 17, 4, 9, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 16, 17, 2, 4, 4, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 3, 3, 20, 2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 18, 2, 18, 4, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2)
                );
    constant threshold_int : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((576, 320, 2112, 1856, 448, 1728, 960, 0, 0, 0, 0, 0, 0, 0, 0),
                (576, 320, 1984, 1728, 320, 1088, 960, 0, 0, 0, 0, 0, 0, 0, 0),
                (576, 320, 2112, 704, 448, 1088, 2368, 0, 0, 0, 0, 0, 0, 0, 0),
                (320, 1984, 576, 576, 576, 576, 1856, 0, 0, 0, 0, 0, 0, 0, 0),
                (448, 1856, 704, 576, 576, 4416, 1984, 0, 0, 0, 0, 0, 0, 0, 0),
                (320, 1728, 576, 576, 960, 1688000, 1728, 0, 0, 0, 0, 0, 0, 0, 0),
                (576, 192, 1984, 1600, 320, 1088, 2368, 0, 0, 0, 0, 0, 0, 0, 0),
                (448, 1600, 704, 576, 704, 576, 1984, 0, 0, 0, 0, 0, 0, 0, 0),
                (576, 704, 1984, 1622976, 192, 960, 2240, 0, 0, 0, 0, 0, 0, 0, 0),
                (320, 1472, 704, 576, 704, 514560, 1984, 0, 0, 0, 0, 0, 0, 0, 0),
                (448, 1600, 576, 576, 832, 1472, 4928, 0, 0, 0, 0, 0, 0, 0, 0),
                (576, 3392, 1856, 192, 704, 1088, 960, 0, 0, 0, 0, 0, 0, 0, 0),
                (1472, 576, 704, 490432, 960, 1620928, 960, 0, 0, 0, 0, 0, 0, 0, 0),
                (320, 1344, 576, 576, 576, 1344, 5440, 0, 0, 0, 0, 0, 0, 0, 0),
                (832, 960, 704, 448, 1837504, 2279936, 960, 0, 0, 0, 0, 0, 0, 0, 0),
                (192, 1216, 704, 960, 1547200, 469952, 2240, 0, 0, 0, 0, 0, 0, 0, 0),
                (1344, 576, 192, 64, 960, 960, 704, 0, 0, 0, 0, 0, 0, 0, 0),
                (576, 2752, 1088, 64, 69312, 960, 2240, 0, 0, 0, 0, 0, 0, 0, 0),
                (1216, 448, 704, 82304, 576, 192, 2368, 0, 0, 0, 0, 0, 0, 0, 0),
                (448, 1344, 576, 576, -71232, 704, 4672, 0, 0, 0, 0, 0, 0, 0, 0),
                (832, 832, 192, 576, 1694656, 960, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (192, 960, 576, 960, 2112, 79360, 4928, 0, 0, 0, 0, 0, 0, 0, 0),
                (704, -74112, 1216, 576, 63104, 2368, 2496, 0, 0, 0, 0, 0, 0, 0, 0),
                (1088, 576, 704, 64, 576, 192, 1216, 0, 0, 0, 0, 0, 0, 0, 0),
                (832, 1344, 576, -86144, 64, 576, 0, 0, 0, 0, 0, 0, 0, -256, -256),
                (192, 1088, 576, 704, -85632, 1620928, 4672, 0, 0, 0, 0, 0, 0, 0, 0),
                (1088, 576, 192, 704, 576, 90432, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (832, 79360, 576, -61632, 576, 64, 704, 0, 0, 0, 0, 0, 0, 0, 0),
                (960, 79872, 704, 448, 576, 476608, 1088, 0, 0, 0, 0, 0, 0, 0, 0),
                (1984, 81792, 448, -72704, 576, 960, 576, 0, 0, 0, 0, 0, 0, 0, 0),
                (576, 1472, 4672, 832, 64, 644608, -43904, 0, 0, 0, 0, 0, 0, 0, 0),
                (704, 432064, 960, 64, 2112, 960, 3520, 0, 0, 0, 0, 0, 0, 0, 0),
                (64, 1205696, 64, 64, 64, 576, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (960, 64, -85632, 1120192, 64, 576, 50112, 0, 0, 0, 0, 0, 0, 0, 0),
                (2276800, 64, 960, 1166784, 64, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (1088, 576, -46720, 704, 3008, 576, 49152, 0, 0, 0, 0, 0, 0, 0, 0),
                (1472, 576, 320, 2234304, 4672, 0, 64, 0, 0, 0, 0, 0, 0, -256, -256),
                (832, 64, 3904, 64, 64, 576, 704, 0, 0, 0, 0, 0, 0, 0, 0),
                (832, -55872, 91904, 0, 75072, -57792, 576, 0, 0, 0, 0, 0, 0, -256, -256),
                (960, 448, 1601472, 64, 74624, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (64, 64, 2279872, 64, 704, 64, 960, 0, 0, 0, 0, 0, 0, 0, 0),
                (960, 1907136, 704, 64, 64, 5952, 3776, 0, 0, 0, 0, 0, 0, 0, 0),
                (1344, 576, 320, 64, 2624, 576, 1077184, 0, 0, 0, 0, 0, 0, 0, 0),
                (-85632, 576, 78912, 320, 192, 704, 704, 0, 0, 0, 0, 0, 0, 0, 0),
                (1600, 576, 1050560, 64, 4672, 0, 1088, 0, 0, 0, 0, 0, 0, -256, -256),
                (832, 304576, 1160128, 576, 767424, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (64, 64, -43904, 64, 704, 576, 42432, 0, 0, 0, 0, 0, 0, 0, 0),
                (99072, 1088, 1216, -98560, 832, 576, 0, 0, 0, 0, 0, 0, 0, -256, -256),
                (1088, 576, 1104832, 496576, 4672, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (1600, 576, 3392, 704, 5568, 1344, 0, 0, 0, 0, 0, 0, 0, -256, -256),
                (704, 1539520, 64, 64, 64, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (64, 64, 1160640, 64, 64, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (1472, 960, 192, -90880, 704, 0, 4672, 0, 0, 0, 0, 0, 0, -256, -256),
                (90880, -36224, 576, -106240, 1088, 320, 0, 0, 0, 0, 0, 0, 0, -256, -256),
                (576, 64, 576, 0, 64, 1600, 4416, 0, 0, 0, 0, 0, 0, -256, -256),
                (46720, -36224, 576, -106240, 64, 320, 4288, 0, 0, 0, 0, 0, 0, 0, 0),
                (5952, 64, 576, 64, 1159104, 320, 960, 0, 0, 0, 0, 0, 0, 0, 0),
                (1344, 576, 448, 64, 1088, 192, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (576, 64, 99072, 0, 64, 832, 576, 0, 0, 0, 0, 0, 0, -256, -256),
                (832, 192, 1088960, 64, 312256, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (5824, 576, 576, 64, 1216, 320, 960, 0, 0, 0, 0, 0, 0, 0, 0),
                (576, 64, 5440, 64, 1582528, 704, 192, 0, 0, 0, 0, 0, 0, 0, 0),
                (704, 1072576, 64, 64, 64, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (99072, 192, 1216, 64, 1008576, 0, 0, 0, 0, 0, 0, -256, -256, -256, -256),
                (5952, 1088, 576, -85632, 832, 1344, -5952, 0, 0, 0, 0, 0, 0, 0, 0),
                (40064, -36224, 576, 576, 576, 320, 3392, 0, 0, 0, 0, 0, 0, 0, 0),
                (1600, 576, 3392, 576, 4416, 1344, 0, 0, 0, 0, 0, 0, 0, -256, -256),
                (1088, 192, 3648, 64, 1077184, 1088, 704, 0, 0, 0, 0, 0, 0, 0, 0),
                (303040, 64, 192, 576, 1088, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (64, 64, 2270144, 737216, 3904, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (1600, 40064, 3392, -46720, 576, 580992, 2624, 0, 0, 0, 0, 0, 0, 0, 0),
                (576, 0, 320, 1023936, 704, 0, 0, 0, 0, -256, -256, -256, -256, -256, -256),
                (378304, 64, 192, 64, 704, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (64, 1088, 2279872, 576, 0, 64, 64, 0, 0, 0, 0, 0, 0, -256, -256),
                (1161152, 64, 64, 64, 64, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (1088, 704, 1213376, 3904, 4672, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (5952, -106240, 576, 704, 64, 1344, 960, 0, 0, 0, 0, 0, 0, 0, 0),
                (704, 105344, 0, 1216, 832, 0, 0, 0, 0, -256, -256, -256, -256, -256, -256),
                (1600, 576, 821184, -59264, 320, 0, 3392, 0, 0, 0, 0, 0, 0, -256, -256),
                (45504, 704, 1216, 64, 2752, 704, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (81792, 832, 704, 192, 64, 2469888, 0, 0, 0, 0, 0, 0, 0, -256, -256),
                (-106240, 320, 960, 576, 0, 960, 832, 0, 0, 0, 0, 0, 0, -256, -256),
                (5824, 1088, 576, 704, 576, -73152, 960, 0, 0, 0, 0, 0, 0, 0, 0),
                (1243584, 64, 64, 64, 320, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (295872, 64, 762304, 576, 448, 1216, 1006016, 0, 0, 0, 0, 0, 0, 0, 0),
                (64, 1646016, 1455552, 64, 64, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (64, 64, 516032, 1014720, 64, 704, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (704, 320, 0, 320, 704, 0, 0, 0, 0, -256, -256, -256, -256, -256, -256),
                (6080, 64, 576, 1088, 64, 0, 0, 0, 0, 0, 0, -256, -256, -256, -256),
                (378304, 64, 762304, 1088, 64, 1216, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (704, 64, 0, 192, 1455552, 0, 0, 0, 0, -256, -256, -256, -256, -256, -256),
                (40064, -36224, 704, 576, 576, 576, 3008, 0, 0, 0, 0, 0, 0, 0, 0),
                (2624, 448, 1856, 576, 448, 0, 64, 0, 0, 0, 0, 0, 0, -256, -256),
                (5952, 320, 576, 320, 576, 320, 0, 0, 0, 0, 0, 0, 0, -256, -256),
                (110080, 1600, 0, 64, 64, 0, 0, 0, 0, -256, -256, -256, -256, -256, -256),
                (-108160, 192, 64, 0, 0, 1088, 192, 0, 0, 0, 0, -256, -256, -256, -256),
                (64, 1728, 704, 1216, 722880, 576, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (64, 3904, 295872, 960, 576, 576, 1728, 0, 0, 0, 0, 0, 0, 0, 0),
                (105792, 832, 832, 192, 704, 0, 0, 0, 0, 0, 0, -256, -256, -256, -256),
                (6080, 39552, 1216, -36224, 576, 0, 0, 0, 0, 0, 0, -256, -256, -256, -256)
                );
    constant children_left : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 13, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 13, 7, 9, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 13, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 13, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 13, 7, 9, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 13, 7, 9, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 9, 3, 5, 7, -1, -1, -1, -1, 11, 13, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 13, 9, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 9, 5, 7, -1, -1, -1, -1, 11, 13, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 13, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 13, 9, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 9, 5, 7, -1, -1, -1, -1, 11, 13, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 9, 5, 7, -1, -1, -1, -1, 11, 13, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 13, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 9, 5, 7, -1, -1, -1, -1, 11, 13, -1, -1, -1, -1),
                (1, 3, 5, 11, 13, 7, 9, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1)
                );
    constant children_right : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 14, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 14, 8, 10, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 14, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 14, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 14, 8, 10, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 14, 8, 10, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 10, 4, 6, 8, -1, -1, -1, -1, 12, 14, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 14, 10, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 10, 6, 8, -1, -1, -1, -1, 12, 14, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 14, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 14, 10, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 10, 6, 8, -1, -1, -1, -1, 12, 14, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 10, 6, 8, -1, -1, -1, -1, 12, 14, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 14, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 10, 6, 8, -1, -1, -1, -1, 12, 14, -1, -1, -1, -1),
                (2, 4, 6, 12, 14, 8, 10, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1)
                );
    constant value_int : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((0, 0, 0, 0, 0, 0, 0, 20, -12, -17, -31, 34, 24, 8, -18),
                (0, 0, 0, 0, 0, 0, 0, 19, -7, -26, -7, 30, 23, 11, -15),
                (0, 0, 0, 0, 0, 0, 0, 14, -13, -11, -24, 27, 19, 6, -15),
                (0, 0, 0, 0, 0, 0, 0, 12, 24, -13, 8, -11, -23, 19, -11),
                (0, 0, 0, 0, 0, 0, 0, 10, 23, -11, 8, -22, -11, 19, -7),
                (0, 0, 0, 0, 0, 0, 0, 12, 22, 9, -12, -18, 1, 18, -7),
                (0, 0, 0, 0, 0, 0, 0, 17, 0, -15, 5, 21, 13, 6, -13),
                (0, 0, 0, 0, 0, 0, 0, 12, 20, -2, 14, -11, -21, 16, -5),
                (0, 0, 0, 0, 0, 0, 0, -2, 18, -6, -18, 20, 13, 7, -8),
                (0, 0, 0, 0, 0, 0, 0, 13, 19, 1, 13, -17, -5, 16, 0),
                (0, 0, 0, 0, 0, 0, 0, 9, 18, 6, -8, 5, -11, -19, -7),
                (0, 0, 0, 0, 0, 0, 0, -3, -15, 9, -8, 17, 8, 5, -10),
                (0, 0, 0, 0, 0, 0, 0, -4, 11, 18, 10, -8, 7, 12, -8),
                (0, 0, 0, 0, 0, 0, 0, 12, 17, -2, 8, 9, -6, -17, -2),
                (0, 0, 0, 0, 0, 0, 0, 15, -2, 0, 14, -14, 0, 8, -7),
                (0, 0, 0, 0, 0, 0, 0, 14, -7, 1, 9, -14, -2, 12, -6),
                (0, 0, 0, 0, 0, 0, 0, 8, -14, 16, 6, 7, -6, -8, 5),
                (0, 0, 0, 0, 0, 0, 0, -9, -19, 4, -17, 14, -10, 4, -6),
                (0, 0, 0, 0, 0, 0, 0, 14, -8, -5, 14, 8, -6, 9, -8),
                (0, 0, 0, 0, 0, 0, 0, 6, 14, -14, 3, 0, -10, -16, -6),
                (0, 0, 0, 0, 0, 0, 0, 5, 14, 0, 11, 1, -5, -13, -5),
                (0, 0, 0, 0, 0, 0, 0, 12, -11, 5, -2, 0, -17, -15, -4),
                (0, 0, 0, 0, 0, 0, 0, -18, -7, 2, -13, 16, 9, 3, -11),
                (0, 0, 0, 0, 0, 0, 0, 9, -9, 15, 9, 6, -4, 9, 2),
                (0, 0, 0, 0, 0, 0, -15, -17, 6, -7, 1, -8, -3, -15, -15),
                (0, 0, 0, 0, 0, 0, 0, 13, 1, -14, 4, -3, 6, -14, -4),
                (0, 0, 0, 0, 0, 0, 0, 13, 0, 14, 7, 3, -17, -6, 1),
                (0, 0, 0, 0, 0, 0, 0, -9, 4, -18, 0, 0, -6, -14, 0),
                (0, 0, 0, 0, 0, 0, 0, 12, 3, -13, 2, -8, 0, 9, 2),
                (0, 0, 0, 0, 0, 0, 0, -10, 4, -17, 0, -8, -1, -7, -13),
                (0, 0, 0, 0, 0, 0, 0, 4, -3, -9, -2, -15, -10, -11, 0),
                (0, 0, 0, 0, 0, 0, 0, 8, -11, -5, 3, 11, -11, 5, -3),
                (0, 0, 0, 0, 0, 0, 0, 6, -23, -14, 5, -14, 0, 6, -4),
                (0, 0, 0, 0, 0, 0, 0, -10, 9, -6, 13, -16, -2, 1, -6),
                (0, 0, 0, 0, 0, 0, 0, -18, 0, -10, 4, 17, 7, 5, -5),
                (0, 0, 0, 0, 0, 0, 0, 10, 0, 15, 8, -9, -1, 1, -5),
                (0, 0, 0, 0, 0, -18, 0, 1, 8, -11, -1, -7, -1, -18, -18),
                (0, 0, 0, 0, 0, 0, 0, -15, 4, -9, 5, -8, 0, -8, 0),
                (0, 0, 0, 0, 0, 0, 0, 10, 0, -6, 1, -14, 0, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, 5, 10, 3, -13, -9, 1, -14, 5),
                (0, 0, 0, 0, 0, 0, 0, 6, 17, 8, 2, -4, 1, 8, -2),
                (0, 0, 0, 0, 0, 0, 0, -5, 2, -12, 7, -16, 0, -6, 1),
                (0, 0, 0, 0, 0, 0, 0, 1, -12, 10, 1, -19, -8, -4, 1),
                (0, 0, 0, 0, 0, 0, 0, -14, -3, 2, -5, 2, -2, -10, 4),
                (0, 0, 0, 0, 0, -12, 0, 4, 0, -9, -1, -10, -2, -12, -12),
                (0, 0, 0, 0, 0, 0, 0, -3, 8, 11, 6, -14, 0, -11, 4),
                (0, 0, 0, 0, 0, 0, 0, 4, 15, 7, 2, -7, -1, 1, -4),
                (0, 0, 0, 0, 0, 0, 0, -12, 1, -16, -4, 0, -14, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, -3, 5, 12, 4, -13, 0, -9, 3),
                (0, 0, 0, 0, 0, 0, -14, 8, 0, -8, 4, -9, -2, -14, -14),
                (0, 0, 0, 0, 0, 0, 0, -6, 2, 9, -1, -8, -2, 8, -1),
                (0, 0, 0, 0, 0, 0, 0, 4, 14, 3, -1, -11, 0, -8, 3),
                (0, 0, 0, 0, 0, -18, 0, -9, 1, -12, -2, -2, -10, -18, -18),
                (0, 0, 0, 0, 0, 0, 0, -12, -2, 1, -5, -13, 0, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, 4, 13, 0, -6, -8, 0, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, -11, -2, 4, 0, -7, 0, 6, -2),
                (0, 0, 0, 0, 0, 0, 0, 7, 1, -2, 1, 9, 20, -6, 4),
                (0, 0, 0, 0, 0, 0, 0, 1, -10, 12, 1, -18, -8, 0, -5),
                (0, 0, 0, 0, 0, 0, 0, 4, 13, 0, -2, -10, 0, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, 0, 10, -2, 4, -10, 0, -7, 2),
                (0, 0, 0, 0, 0, 0, 0, 0, -10, 5, -3, 7, 14, -5, 4),
                (0, 0, 0, 0, 0, 0, 0, -1, 10, -1, 2, -5, -14, 8, -2),
                (0, 0, 0, 0, 0, 0, 0, -9, 1, -5, 4, -7, -1, 7, 0),
                (0, 0, 0, 0, 0, -9, 0, -7, 2, -8, 0, -9, -9, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, -6, 0, -14, -2, 11, 0, 0, -6),
                (0, 0, 0, 0, 0, 0, 0, -3, 0, 2, 0, -5, 0, 6, -2),
                (0, 0, 0, 0, 0, 0, -11, 7, 0, -6, 0, -6, 0, -11, -11),
                (0, 0, 0, 0, 0, 0, 0, -7, 2, -6, 1, -12, -5, -10, 2),
                (0, 0, 0, 0, 0, 0, 0, -14, 2, 3, -3, 1, 13, -8, 0),
                (0, 0, 0, 0, 0, 0, 0, 11, 2, 3, -1, -4, 0, 10, 0),
                (0, 0, 0, 0, 0, 0, 0, -2, 1, -3, 2, -8, -1, -12, 0),
                (0, 6, 0, 0, 0, -6, 2, 1, -1, 6, 6, 6, 6, 6, 6),
                (0, 0, 0, 0, 0, 0, 0, 32, 2, -6, 2, 5, -2, -7, 0),
                (0, 0, 0, 0, -20, 0, 0, -3, 15, -2, 1, 9, 0, -20, -20),
                (0, 0, 0, 0, 0, 0, 0, 22, -11, 1, -6, 8, -7, -9, 1),
                (0, 0, 0, 0, 0, 0, 0, -2, 2, 10, 2, -7, 0, 5, -1),
                (0, 0, 0, 0, 0, 0, 0, -10, 0, 2, 0, 10, 0, -4, 4),
                (0, 0, -11, 0, 0, 0, -5, -10, 0, -11, -11, -11, -11, -11, -11),
                (0, 0, 0, 0, 0, -6, 0, 0, 7, -2, 0, -1, -8, -6, -6),
                (0, 0, 0, 0, 0, 0, 0, 1, -9, 6, -4, 12, 1, -9, 0),
                (0, 0, 0, 0, 0, 0, 2, 7, 1, 1, 0, -5, 4, 2, 2),
                (0, 0, 0, 0, 0, 0, 0, -12, 0, 2, 0, -9, 0, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, -1, 1, -2, -12, 0, 7, -4, 3),
                (0, 0, 0, 0, 0, 0, 0, -5, 1, -13, -1, 0, -13, -4, 3),
                (0, 0, 0, 0, 0, 0, 0, -12, 2, -5, 1, 4, -1, -3, 1),
                (0, 0, 0, 0, 0, 0, 0, 0, -3, 13, 1, 18, 3, -13, -1),
                (0, 0, 0, 0, 0, 0, 0, -9, 1, 27, 3, -4, 2, 1, -5),
                (0, 0, -10, 0, 0, -4, 4, 1, -1, -10, -10, -10, -10, -10, -10),
                (0, 0, 0, 0, 0, 15, 0, 7, -18, 0, -1, 15, 15, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, -2, -14, 5, -1, 4, 0, 0, -8),
                (0, 0, -10, 0, 0, 6, 0, 9, -2, -10, -10, -10, -10, -10, -10),
                (0, 0, 0, 0, 0, 0, 0, -2, 0, 2, 0, -3, 1, 5, -2),
                (0, 0, 0, 0, 0, -10, 0, 1, -4, 1, -2, 5, -5, -10, -10),
                (0, 0, 0, 0, 0, 0, -1, -4, 2, 0, -4, 4, 11, -1, -1),
                (0, 0, -8, 0, 0, -1, 1, -2, -6, -8, -8, -8, -8, -8, -8),
                (0, 0, 0, 0, -10, 0, 0, 1, -1, 10, 0, 0, 0, -10, -10),
                (0, 0, 0, 0, 0, 0, 0, -11, -1, 8, 1, -2, 5, 0, -2),
                (0, 0, 0, 0, 0, 0, 0, 7, 2, 4, -4, -4, 1, -1, 1),
                (0, 0, 0, 0, 0, -8, 0, 2, 0, -5, 0, -8, -8, 0, 0),
                (0, 0, 0, 0, 0, 13, 0, -1, 1, -2, 0, 13, 13, 0, 0)
                );
    constant parent : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 6, 6, 5, 5),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 4, 4, 5, 5, 6, 6, 3, 3),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 6, 6, 5, 5),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 6, 6, 5, 5),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 4, 4, 5, 5, 6, 6, 3, 3),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 4, 4, 5, 5, 6, 6, 3, 3),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 2, 2, 3, 3, 4, 4, 1, 1, 9, 9, 10, 10),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 5, 5, 6, 6, 4, 4),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 3, 3, 4, 4, 2, 2, 9, 9, 10, 10),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 6, 6, 5, 5),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 5, 5, 6, 6, 4, 4),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 3, 3, 4, 4, 2, 2, 9, 9, 10, 10),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 3, 3, 4, 4, 2, 2, 9, 9, 10, 10),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 6, 6, 5, 5),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 3, 3, 4, 4, 2, 2, 9, 9, 10, 10),
                (-1, 0, 0, 1, 1, 2, 2, 5, 5, 6, 6, 3, 3, 4, 4),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6)
                );
    constant depth : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 3, 3, 3, 3, 2, 2, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 3, 3, 3, 3, 2, 2, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 3, 3, 3, 3, 2, 2, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 3, 3, 3, 3, 2, 2, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 3, 3, 3, 3, 2, 2, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3)
                );
    constant iLeaf : intArray2D(nTrees-1 downto 0)(nLeaves-1 downto 0) := ((7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (5, 6, 7, 8, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (5, 6, 7, 8, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (5, 6, 7, 8, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (5, 6, 7, 8, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (5, 6, 7, 8, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14)
                );
    constant value : tyArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := to_tyArray2D(value_int);
      constant threshold : txArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := to_txArray2D(threshold_int);
end Arrays0;