LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;


use work.ipbus.all;
use work.emp_data_types.all;
use work.emp_project_decl.all;

use work.emp_device_decl.all;
use work.emp_ttc_decl.all;

--library GBDT;
use work.Constants.all;
use work.Types.all;


entity NNWrapper is
  port (
    ap_clk : in std_logic;
    LinksIn : in ldata(4 * N_REGION - 1 downto 0) := ( others => LWORD_NULL );
    LinksOut : out ldata(4 * N_REGION - 1 downto 0) := ( others => LWORD_NULL );
    ap_rst : in std_logic;
    
    ap_done : out std_logic;
    ap_idle : out std_logic;
    ap_ready : out std_logic
    
  );
end entity NNWrapper;

architecture rtl of NNWrapper is
  signal input_1_V_ap_vld : STD_LOGIC := '0';
  signal input_1_V : STD_LOGIC_VECTOR (NN_bit_width*nFeatures -1 downto 0);
  signal layer13_out_0_V : STD_LOGIC_VECTOR (NN_bit_width -1 downto 0);
  signal layer13_out_0_V_ap_vld : STD_LOGIC := '0';

  signal X : txArray(0 to nFeatures - 1) := (others => to_tx(0));
  signal X_vld : boolean := false;

  signal ap_start : std_logic := '0';

  signal const_size_in_1 : STD_LOGIC_VECTOR (NN_bit_width -1 downto 0);
  signal const_size_in_1_ap_vld : std_logic := '0';
  signal const_size_out_1 : STD_LOGIC_VECTOR (NN_bit_width -1 downto 0);
  signal const_size_out_1_ap_vld : std_logic := '0';

begin

    Input : entity work.FeatureTransform
    port map(ap_clk, X, X_vld,LinksIn);

    UIN : entity work.RunningInput
    port map(ap_clk, input_1_V_ap_vld, input_1_V,X,X_vld,ap_start);

    UUT : entity work.myproject
    port map( ap_clk,
              ap_rst,
              ap_start,
              ap_done,
              ap_idle,
              ap_ready,
              input_1_V_ap_vld,
              input_1_V,
              layer13_out_0_V,
              layer13_out_0_V_ap_vld,
              const_size_in_1,
              const_size_in_1_ap_vld,
              const_size_out_1,
              const_size_out_1_ap_vld);

    Output : entity work.RunningOutput
    port map(ap_clk, layer13_out_0_V,layer13_out_0_V_ap_vld,LinksOut);

end architecture rtl;
