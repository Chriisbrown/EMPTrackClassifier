library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_misc.all;
  use ieee.numeric_std.all;

  use work.Constants.all;
  use work.Types.all;
  package Arrays0 is

    constant initPredict : ty := to_ty(0);
    constant feature : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((4, 1, 0, 0, 1, 0, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 1, 0, 0, 19, 2, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 1, 0, 3, 1, 2, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 4, 4, 4, 3, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 4, 4, 4, 16, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 4, 4, 3, 17, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 1, 0, 0, 19, 2, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 4, 4, 4, 1, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 3, 0, 17, 1, 2, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 4, 4, 4, 17, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 1, 4, 3, 0, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 16, 0, 1, 3, 2, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 4, 4, 17, 2, 17, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 1, 4, 4, 0, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 2, 4, 1, 17, 17, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 2, 4, 3, 17, 17, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 4, 1, 10, 2, 3, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 16, 2, 10, 18, 3, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 1, 4, 18, 4, 20, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 1, 4, 18, 3, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 2, 1, 4, 17, 3, 12, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 2, 1, 3, 0, 18, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 18, 2, 4, 18, 16, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 4, 4, 10, 2, 20, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 2, 1, 18, 7, 4, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 1, 2, 18, 17, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 4, 1, 0, 2, 18, 12, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 18, 1, 18, 4, 5, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 18, 4, 1, 4, 17, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 18, 1, 18, 4, 16, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 2, 16, 3, 7, 17, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 17, 2, 5, 16, 3, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (7, 17, 6, 5, 12, 20, 13, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 7, 18, 17, 6, 4, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 7, 3, 17, 6, 14, 14, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 4, 18, 0, 16, 4, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 1, 16, 17, 16, -2, 12, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 7, 16, 13, 6, 20, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 18, 18, -2, 18, 18, 20, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 2, 17, 7, 18, 7, 12, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 5, 17, 8, 2, 7, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 17, 2, 7, 13, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 20, 16, 10, 16, 20, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 4, 18, 19, 1, 3, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 1, 17, 5, 16, -2, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 17, 17, 4, 17, 7, 12, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 5, 18, 8, 2, 4, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 3, 3, 18, 2, 16, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 20, 17, 17, 16, 7, 12, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 1, 16, 0, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2, -2)
                );
    constant threshold_int : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((576, 2, 2112, 1856, 4, 1728, 8, 0, 0, 0, 0, 0, 0, 0, 0),
                (576, 2, 1984, 1728, 320, 8, 8, 0, 0, 0, 0, 0, 0, 0, 0),
                (576, 2, 2112, 6, 4, 8, 2368, 0, 0, 0, 0, 0, 0, 0, 0),
                (2, 1984, 576, 576, 576, 4, 1856, 0, 0, 0, 0, 0, 0, 0, 0),
                (4, 1856, 704, 576, 576, 34, 1984, 0, 0, 0, 0, 0, 0, 0, 0),
                (2, 1728, 576, 576, 8, 13188, 1728, 0, 0, 0, 0, 0, 0, 0, 0),
                (576, 2, 1984, 1600, 320, 8, 2368, 0, 0, 0, 0, 0, 0, 0, 0),
                (4, 1600, 704, 576, 704, 4, 1984, 0, 0, 0, 0, 0, 0, 0, 0),
                (576, 6, 1984, 12680, 2, 8, 2240, 0, 0, 0, 0, 0, 0, 0, 0),
                (2, 1472, 704, 576, 704, 4020, 1984, 0, 0, 0, 0, 0, 0, 0, 0),
                (4, 1600, 4, 576, 6, 1472, 38, 0, 0, 0, 0, 0, 0, 0, 0),
                (576, 26, 1856, 2, 6, 8, 8, 0, 0, 0, 0, 0, 0, 0, 0),
                (1472, 576, 704, 3832, 8, 12664, 8, 0, 0, 0, 0, 0, 0, 0, 0),
                (2, 1344, 4, 576, 576, 1344, 42, 0, 0, 0, 0, 0, 0, 0, 0),
                (6, 8, 704, 4, 14356, 17812, 8, 0, 0, 0, 0, 0, 0, 0, 0),
                (2, 10, 704, 8, 12088, 3672, 2240, 0, 0, 0, 0, 0, 0, 0, 0),
                (1344, 576, 2, 64, 8, 8, 704, 0, 0, 0, 0, 0, 0, 0, 0),
                (576, 22, 8, 64, 542, 8, 2240, 0, 0, 0, 0, 0, 0, 0, 0),
                (1216, 4, 704, 643, 576, 192, 2368, 0, 0, 0, 0, 0, 0, 0, 0),
                (4, 1344, 4, 576, -556, 6, 36, 0, 0, 0, 0, 0, 0, 0, 0),
                (6, 6, 2, 576, 13240, 8, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (2, 8, 4, 8, 2112, 620, 38, 0, 0, 0, 0, 0, 0, 0, 0),
                (704, -579, 10, 576, 493, 18, 2496, 0, 0, 0, 0, 0, 0, 0, 0),
                (1088, 576, 704, 64, 4, 192, 10, 0, 0, 0, 0, 0, 0, 0, 0),
                (6, 10, 4, -673, 64, 576, 0, 0, 0, 0, 0, 0, 0, -256, -256),
                (2, 1088, 4, 6, -669, 12664, 36, 0, 0, 0, 0, 0, 0, 0, 0),
                (1088, 576, 2, 704, 4, 706, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (6, 620, 4, -482, 576, 64, 704, 0, 0, 0, 0, 0, 0, 0, 0),
                (960, 624, 704, 4, 576, 3724, 8, 0, 0, 0, 0, 0, 0, 0, 0),
                (1984, 639, 4, -568, 576, 8, 4, 0, 0, 0, 0, 0, 0, 0, 0),
                (4, 12, 36, 6, 64, 5036, -343, 0, 0, 0, 0, 0, 0, 0, 0),
                (704, 3376, 8, 64, 16, 8, 28, 0, 0, 0, 0, 0, 0, 0, 0),
                (64, 9420, 64, 64, 64, 576, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (960, 64, -669, 8752, 64, 576, 392, 0, 0, 0, 0, 0, 0, 0, 0),
                (17788, 64, 8, 9116, 64, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (1088, 576, -365, 704, 24, 576, 384, 0, 0, 0, 0, 0, 0, 0, 0),
                (12, 4, 2, 17456, 36, 0, 64, 0, 0, 0, 0, 0, 0, -256, -256),
                (6, 64, 30, 64, 64, 576, 6, 0, 0, 0, 0, 0, 0, 0, 0),
                (832, -436, 718, 0, 586, -452, 576, 0, 0, 0, 0, 0, 0, -256, -256),
                (960, 4, 12512, 64, 583, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (0, 64, 17812, 64, 6, 64, 8, 0, 0, 0, 0, 0, 0, 0, 0),
                (8, 14900, 6, 64, 64, 46, 30, 0, 0, 0, 0, 0, 0, 0, 0),
                (10, 576, 2, 64, 20, 576, 8416, 0, 0, 0, 0, 0, 0, 0, 0),
                (-669, 576, 616, 320, 2, 6, 704, 0, 0, 0, 0, 0, 0, 0, 0),
                (12, 4, 8208, 64, 36, 0, 8, 0, 0, 0, 0, 0, 0, -256, -256),
                (832, 2380, 9064, 576, 5996, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (0, 64, -343, 64, 6, 576, 332, 0, 0, 0, 0, 0, 0, 0, 0),
                (774, 8, 10, -770, 6, 4, 0, 0, 0, 0, 0, 0, 0, -256, -256),
                (1088, 576, 8632, 3880, 36, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (12, 4, 26, 704, 44, 10, 0, 0, 0, 0, 0, 0, 0, -256, -256)
                );
    constant children_left : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 13, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 13, 7, 9, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 13, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1)
                );
    constant children_right : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 14, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 14, 8, 10, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 14, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1)
                );
    constant value_int : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((0, 0, 0, 0, 0, 0, 0, 20, -12, -17, -31, 34, 24, 8, -18),
                (0, 0, 0, 0, 0, 0, 0, 19, -7, -26, -7, 30, 23, 11, -15),
                (0, 0, 0, 0, 0, 0, 0, 14, -13, -11, -24, 27, 19, 6, -15),
                (0, 0, 0, 0, 0, 0, 0, 12, 24, -13, 8, -11, -23, 19, -11),
                (0, 0, 0, 0, 0, 0, 0, 10, 23, -11, 8, -22, -11, 19, -7),
                (0, 0, 0, 0, 0, 0, 0, 12, 22, 9, -12, -18, 1, 18, -7),
                (0, 0, 0, 0, 0, 0, 0, 17, 0, -15, 5, 21, 13, 6, -13),
                (0, 0, 0, 0, 0, 0, 0, 12, 20, -2, 14, -11, -21, 16, -5),
                (0, 0, 0, 0, 0, 0, 0, -2, 18, -6, -18, 20, 13, 7, -8),
                (0, 0, 0, 0, 0, 0, 0, 13, 19, 1, 13, -17, -5, 16, 0),
                (0, 0, 0, 0, 0, 0, 0, 9, 18, 6, -8, 5, -11, -19, -7),
                (0, 0, 0, 0, 0, 0, 0, -3, -15, 9, -8, 17, 8, 5, -10),
                (0, 0, 0, 0, 0, 0, 0, -4, 11, 18, 10, -8, 7, 12, -8),
                (0, 0, 0, 0, 0, 0, 0, 12, 17, -2, 8, 9, -6, -17, -2),
                (0, 0, 0, 0, 0, 0, 0, 15, -2, 0, 14, -14, 0, 8, -7),
                (0, 0, 0, 0, 0, 0, 0, 14, -7, 1, 9, -14, -2, 12, -6),
                (0, 0, 0, 0, 0, 0, 0, 8, -14, 16, 6, 7, -6, -8, 5),
                (0, 0, 0, 0, 0, 0, 0, -9, -19, 4, -17, 14, -10, 4, -6),
                (0, 0, 0, 0, 0, 0, 0, 14, -8, -5, 14, 8, -6, 9, -8),
                (0, 0, 0, 0, 0, 0, 0, 6, 14, -14, 3, 0, -10, -16, -6),
                (0, 0, 0, 0, 0, 0, 0, 5, 14, 0, 11, 1, -5, -13, -5),
                (0, 0, 0, 0, 0, 0, 0, 12, -11, 5, -2, 0, -17, -15, -4),
                (0, 0, 0, 0, 0, 0, 0, -18, -7, 2, -13, 16, 9, 3, -11),
                (0, 0, 0, 0, 0, 0, 0, 9, -9, 15, 9, 6, -4, 9, 2),
                (0, 0, 0, 0, 0, 0, -15, -17, 6, -7, 1, -8, -3, -15, -15),
                (0, 0, 0, 0, 0, 0, 0, 13, 1, -14, 4, -3, 6, -14, -4),
                (0, 0, 0, 0, 0, 0, 0, 13, 0, 14, 7, 3, -17, -6, 1),
                (0, 0, 0, 0, 0, 0, 0, -9, 4, -18, 0, 0, -6, -14, 0),
                (0, 0, 0, 0, 0, 0, 0, 12, 3, -13, 2, -8, 0, 9, 2),
                (0, 0, 0, 0, 0, 0, 0, -10, 4, -17, 0, -8, -1, -7, -13),
                (0, 0, 0, 0, 0, 0, 0, 4, -3, -9, -2, -15, -10, -11, 0),
                (0, 0, 0, 0, 0, 0, 0, 8, -11, -5, 3, 11, -11, 5, -3),
                (0, 0, 0, 0, 0, 0, 0, 6, -23, -14, 5, -14, 0, 6, -4),
                (0, 0, 0, 0, 0, 0, 0, -10, 9, -6, 13, -16, -2, 1, -6),
                (0, 0, 0, 0, 0, 0, 0, -18, 0, -10, 4, 17, 7, 5, -5),
                (0, 0, 0, 0, 0, 0, 0, 10, 0, 15, 8, -9, -1, 1, -5),
                (0, 0, 0, 0, 0, -18, 0, 1, 8, -11, -1, -7, -1, -18, -18),
                (0, 0, 0, 0, 0, 0, 0, -15, 4, -9, 5, -8, 0, -8, 0),
                (0, 0, 0, 0, 0, 0, 0, 10, 0, -6, 1, -14, 0, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, 5, 10, 3, -13, -9, 1, -14, 5),
                (0, 0, 0, 0, 0, 0, 0, 6, 17, 8, 2, -4, 1, 8, -2),
                (0, 0, 0, 0, 0, 0, 0, -5, 2, -12, 7, -16, 0, -6, 1),
                (0, 0, 0, 0, 0, 0, 0, 1, -12, 10, 1, -19, -8, -4, 1),
                (0, 0, 0, 0, 0, 0, 0, -14, -3, 2, -5, 2, -2, -10, 4),
                (0, 0, 0, 0, 0, -12, 0, 4, 0, -9, -1, -10, -2, -12, -12),
                (0, 0, 0, 0, 0, 0, 0, -3, 8, 11, 6, -14, 0, -11, 4),
                (0, 0, 0, 0, 0, 0, 0, 4, 15, 7, 2, -7, -1, 1, -4),
                (0, 0, 0, 0, 0, 0, 0, -12, 1, -16, -4, 0, -14, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, -3, 5, 12, 4, -13, 0, -9, 3),
                (0, 0, 0, 0, 0, 0, -14, 8, 0, -8, 4, -9, -2, -14, -14)
                );
    constant parent : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 6, 6, 5, 5),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 4, 4, 5, 5, 6, 6, 3, 3),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 6, 6, 5, 5),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6)
                );
    constant depth : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3)
                );
    constant iLeaf : intArray2D(nTrees-1 downto 0)(nLeaves-1 downto 0) := ((7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14)
                );
    constant value : tyArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := to_tyArray2D(value_int);
      constant threshold : txArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := to_txArray2D(threshold_int);
end Arrays0;