library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_misc.all;
  use ieee.numeric_std.all;

  use work.Constants.all;
  use work.Types.all;
  package Arrays0 is

    constant initPredict : ty := to_ty(0);
    constant feature : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((4, 1, 0, 3, 1, 0, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 1, 0, 0, 19, 3, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 4, 0, 3, 1, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 17, 0, 0, 3, 0, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 1, 18, 4, 3, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 3, 3, 18, 1, 0, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 1, 17, 2, 4, 1, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 1, 3, 4, 17, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 0, 4, 4, 5, 5, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 17, 16, 5, 3, 0, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 7, 14, 17, 6, 15, 12, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 16, 18, 16, 1, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 3, 4, 2, 12, 1, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 7, 13, 5, 13, 15, 12, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 16, 2, 17, 16, 19, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 7, 16, 12, 6, 20, 19, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 5, 16, 8, 16, 3, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 18, 16, 1, 17, 16, 10, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 0, 2, 1, 17, 20, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (19, 11, 17, 0, 16, 7, 12, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 15, 16, 17, 13, 17, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (7, 13, 13, 10, 12, 17, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 17, 8, 7, 14, 10, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 3, 4, 16, 16, 0, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 16, 2, 4, 2, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 0, 18, 4, 3, 4, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 17, 10, 4, 17, 3, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (10, 4, 4, 16, 16, 7, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 1, 17, 5, 18, 11, 19, -2, -2, -2, -2, -2, -2, -2, -2),
                (7, 17, 4, 5, 16, 10, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 17, 4, 5, 2, 1, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 16, 16, 4, 16, 9, 10, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 16, 18, 17, 4, 4, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 17, 19, 4, 17, 14, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 20, 14, 11, 5, 15, 19, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 16, 17, 0, 17, 16, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 17, 6, 17, 2, 19, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 7, 17, 4, 2, 15, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 1, 0, 1, 3, 1, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 3, 0, 5, 1, 3, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 17, 10, 6, 1, 3, 7, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 0, 18, 0, 17, 1, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 2, 16, 17, 5, 3, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (20, 4, 19, 12, 2, 17, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 17, 0, -2, 0, 17, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 16, 4, 4, 12, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 16, 16, 20, 2, 0, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 17, 2, 5, 2, 20, 20, -2, -2, -2, -2, -2, -2, -2, -2),
                (8, 16, 3, 4, 0, 9, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 18, 0, 0, 0, 2, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 16, 16, 4, 17, 17, 20, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 16, 1, 3, 0, 4, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 4, 18, 15, 2, 0, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 5, 3, 16, 16, 16, 6, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 18, 18, 18, 20, 4, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 20, 14, 11, 17, 15, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 3, 14, 3, 17, 6, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 0, 16, 2, 3, 20, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (5, 17, 1, 2, 17, 15, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 5, 3, 17, 16, 10, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 4, 4, 2, 0, 0, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 17, 16, 7, 14, 0, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 20, 2, 17, 0, 7, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 4, 18, 16, 16, 16, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 14, 1, 0, 2, 4, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 10, 17, 9, 4, 4, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 0, 17, 3, 16, 3, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 3, 1, 1, 0, 1, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 3, 17, 3, 1, 16, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 16, 18, 1, 18, 1, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 18, 18, 1, 0, 1, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 2, 17, 0, 17, 18, 19, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 20, 2, 0, 17, 19, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (5, 1, 1, 17, 7, 1, 7, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 16, 4, 2, 3, 16, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 2, 20, 16, 16, 0, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 0, 3, 16, -2, 4, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 17, 4, 18, 17, 6, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 16, 1, 16, 1, 16, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 18, 0, 10, 2, 16, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 2, 16, 10, 3, 9, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 3, 17, 16, 3, 0, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 3, 20, 6, 19, 10, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (19, 17, 12, 13, 15, 15, 15, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 20, 15, 4, 0, 2, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 4, 3, 0, 18, 2, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 1, 1, 3, 1, 17, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 0, 0, 16, 16, 1, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 0, 4, 17, 20, 15, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 17, 14, 2, 14, 15, 19, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 3, 1, 3, 17, 2, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 1, 3, 1, 10, 1, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 1, 0, 16, 0, 2, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 14, 0, 6, 16, 2, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 3, 3, 1, 1, 4, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 16, 16, 2, 0, 0, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 2, 18, 18, 16, 0, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 17, 0, 17, 17, 4, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 15, 16, 5, 12, 4, 7, -2, -2, -2, -2, -2, -2, -2, -2),
                (8, 10, 3, 17, 2, 9, 6, -2, -2, -2, -2, -2, -2, -2, -2)
                );
    constant threshold_int : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((576, 60, 428, 178, 117, 333, 258, 0, 0, 0, 0, 0, 0, 0, 0),
                (576, 37, 470, 380, 320, 289, 96, 0, 0, 0, 0, 0, 0, 0, 0),
                (105, 354, 704, 268, 236, 168, 601, 0, 0, 0, 0, 0, 0, 0, 0),
                (576, 396, 578, 208, 206, 309, 213, 0, 0, 0, 0, 0, 0, 0, 0),
                (129, 535, 183, 1271, 704, 164, 302014, 0, 0, 0, 0, 0, 0, 0, 0),
                (704, 210, 307, 964, -7, 757, 316, 0, 0, 0, 0, 0, 0, 0, 0),
                (289, 194, 462, 71, 576, 12, 279, 0, 0, 0, 0, 0, 0, 0, 0),
                (144, 721, 212, 270, 576, 114, 301421, 0, 0, 0, 0, 0, 0, 0, 0),
                (1084, 234, 576, 576, 64, 64, 337, 0, 0, 0, 0, 0, 0, 0, 0),
                (704, 124, 172001, 64, 149, 521, 158, 0, 0, 0, 0, 0, 0, 0, 0),
                (546, 64, 64, 289, 64, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (198, 758, 284429, 1534, 27004, 234, 91, 0, 0, 0, 0, 0, 0, 0, 0),
                (656, 318, 704, 9, 64, -39, 222649, 0, 0, 0, 0, 0, 0, 0, 0),
                (386, 64, 64, 64, 64, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (238, 141, 365078, -92, 262, 264242, 320, 0, 0, 0, 0, 0, 0, 0, 0),
                (304, 64, 196502, 64, 64, 576, 576, 0, 0, 0, 0, 0, 0, 0, 0),
                (-86, 64, 372718, 64, 230586, 109, 576, 0, 0, 0, 0, 0, 0, 0, 0),
                (674, 1661, 27498, 253, 617, 10439, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (2964, 292, -78, 61, 4, 576, 270, 0, 0, 0, 0, 0, 0, 0, 0),
                (192, 64, 248, 396, 135183, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (811, 64, 77290, 376, 64, 580, 209115, 0, 0, 0, 0, 0, 0, 0, 0),
                (64, 64, 64, 64, 64, 249, 704, 0, 0, 0, 0, 0, 0, 0, 0),
                (-41, 246, 64, 64, 64, 64, 217084, 0, 0, 0, 0, 0, 0, 0, 0),
                (369721, 329, 576, 318974, 224032, 609, 288, 0, 0, 0, 0, 0, 0, 0, 0),
                (255, 50089, 458, 576, 98, 40901, 85325, 0, 0, 0, 0, 0, 0, 0, 0),
                (5302, 406, 1414, 576, 163, 576, 576, 0, 0, 0, 0, 0, 0, 0, 0),
                (261, 62, 64, 576, 186, 170, 704, 0, 0, 0, 0, 0, 0, 0, 0),
                (64, 576, 576, 175459, 230849, 64, 121945, 0, 0, 0, 0, 0, 0, 0, 0),
                (832, -145, 321, 64, 1661, 64, 576, 0, 0, 0, 0, 0, 0, 0, 0),
                (64, 297, 576, 64, 112625, 64, 297437, 0, 0, 0, 0, 0, 0, 0, 0),
                (360632, 187, 576, 64, 460, 49, 306, 0, 0, 0, 0, 0, 0, 0, 0),
                (625, 24303, 18771, 576, 212276, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (256, 29210, 731, 70, 576, 576, 576, 0, 0, 0, 0, 0, 0, 0, 0),
                (99, 78, 320, 576, 189, 64, 369, 0, 0, 0, 0, 0, 0, 0, 0),
                (300, 320, 64, 64, 64, 64, 320, 0, 0, 0, 0, 0, 0, 0, 0),
                (252, 5467, 108, 406, 731, 324374, 469, 0, 0, 0, 0, 0, 0, 0, 0),
                (442, 187, 64, 105, 451, 576, 102, 0, 0, 0, 0, 0, 0, 0, 0),
                (314, 64, 355, 704, -117, 64, 106368, 0, 0, 0, 0, 0, 0, 0, 0),
                (374331, 281, 231, 104, 1, 50, 633, 0, 0, 0, 0, 0, 0, 0, 0),
                (-79, 468, -25, 64, -170, -424, 273, 0, 0, 0, 0, 0, 0, 0, 0),
                (177, 145, 64, 64, 28, 165, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (11, 363, 484, 213, 652, 128, 576, 0, 0, 0, 0, 0, 0, 0, 0),
                (193, 798, 333694, 687, 64, 154, 464, 0, 0, 0, 0, 0, 0, 0, 0),
                (64, 576, 576, 64, 511, 314, 532, 0, 0, 0, 0, 0, 0, 0, 0),
                (2964, 13, 832, 0, 450, 187, 2, 0, 0, 0, 0, 0, 0, -256, -256),
                (324, 62273, 576, 576, 64, 139036, 248533, 0, 0, 0, 0, 0, 0, 0, 0),
                (704, 100737, 132483, 576, 355, 418, 219, 0, 0, 0, 0, 0, 0, 0, 0),
                (275, 639, 72, 64, 169, 576, 576, 0, 0, 0, 0, 0, 0, 0, 0),
                (64, 225053, 136, 704, 730, 64, 308, 0, 0, 0, 0, 0, 0, 0, 0),
                (-468, 1106, 875, 23, 368, 873, 877, 0, 0, 0, 0, 0, 0, 0, 0),
                (535, 53085, 23941, 576, 187, 472, 576, 0, 0, 0, 0, 0, 0, 0, 0),
                (-25, 295131, 38, 360, 631, 576, 259236, 0, 0, 0, 0, 0, 0, 0, 0),
                (229, 576, 386, 64, 158, 319, 1519, 0, 0, 0, 0, 0, 0, 0, 0),
                (536, 64, 256, 157017, 114042, 265197, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (445, 1721, 1616, 1016, 192, 704, 541, 0, 0, 0, 0, 0, 0, 0, 0),
                (308, 320, 64, 64, 290, 64, 337, 0, 0, 0, 0, 0, 0, 0, 0),
                (576, 442, 64, 437, 670, 64, -40, 0, 0, 0, 0, 0, 0, 0, 0),
                (6257, 317, 373969, -153, 212, 64, 375484, 0, 0, 0, 0, 0, 0, 0, 0),
                (64, 175, 109, 226, 241, 64, 246, 0, 0, 0, 0, 0, 0, 0, 0),
                (74, 64, 129, 171, 183823, 64, 454, 0, 0, 0, 0, 0, 0, 0, 0),
                (269610, 576, 576, 326, 378, 603, 268, 0, 0, 0, 0, 0, 0, 0, 0),
                (459, 331, 47619, 64, 64, 446, 166, 0, 0, 0, 0, 0, 0, 0, 0),
                (-129, 576, -127, 103, -82, 64, 704, 0, 0, 0, 0, 0, 0, 0, 0),
                (536, 704, 574, 199005, 98037, 58387, 1331, 0, 0, 0, 0, 0, 0, 0, 0),
                (-242, 64, -221, 154, 324, 576, 964, 0, 0, 0, 0, 0, 0, 0, 0),
                (94, 64, 202, 64, 576, 576, 194, 0, 0, 0, 0, 0, 0, 0, 0),
                (1, 589, 734, 320, 43766, 174, 1211, 0, 0, 0, 0, 0, 0, 0, 0),
                (-82, -436, 104, 42, -221, 86, 1234, 0, 0, 0, 0, 0, 0, 0, 0),
                (12, 98, 13, 88, 118, 149509, 14, 0, 0, 0, 0, 0, 0, 0, 0),
                (-303, 312157, 131, 32, 326, 33, 259, 0, 0, 0, 0, 0, 0, 0, 0),
                (180, 1099, 319, 179, 651, 186, 321, 0, 0, 0, 0, 0, 0, 0, 0),
                (281, 713, 266, 682, 628, 71, 448, 0, 0, 0, 0, 0, 0, 0, 0),
                (557, 64, 103, 423, 526, 448, 367152, 0, 0, 0, 0, 0, 0, 0, 0),
                (64, 142, 96, 170, 64, 86, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (361422, 355396, 704, 538, 182, 361916, -91, 0, 0, 0, 0, 0, 0, 0, 0),
                (237765, 461, 576, 18507, 10505, 711, 496, 0, 0, 0, 0, 0, 0, 0, 0),
                (862, 861, 197, 26279, 0, 704, 236, 0, 0, 0, 0, 0, 0, -256, -256),
                (1714, 2, 704, 64, 11, 64, 677, 0, 0, 0, 0, 0, 0, 0, 0),
                (742, 342882, 95, 342684, 128, 346702, 0, 0, 0, 0, 0, 0, 0, -256, -256),
                (1901, 1879, 484, 64, 402, 317031, 139, 0, 0, 0, 0, 0, 0, 0, 0),
                (301, 530, 208917, 64, 258, 64, 370643, 0, 0, 0, 0, 0, 0, 0, 0),
                (134, 187, 159, 203681, 338, 330, 221, 0, 0, 0, 0, 0, 0, 0, 0),
                (189784, 185, 704, 64, 576, 64, 519, 0, 0, 0, 0, 0, 0, 0, 0),
                (320, 452, 64, 64, 64, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (557, 64, 64, 576, 205, 372, 704, 0, 0, 0, 0, 0, 0, 0, 0),
                (375056, 704, 356, 533, 1189, 518, 442, 0, 0, 0, 0, 0, 0, 0, 0),
                (-387, -495, -371, 24, -459, 335, 463, 0, 0, 0, 0, 0, 0, 0, 0),
                (173, 168, 173, 50385, 286108, 74, -54, 0, 0, 0, 0, 0, 0, 0, 0),
                (68958, 316, 576, 131, 576, 64, -25, 0, 0, 0, 0, 0, 0, 0, 0),
                (331, 329, 64, 261, 64, 64, 320, 0, 0, 0, 0, 0, 0, 0, 0),
                (-153, -100, -152, -101, 537, 140, -127, 0, 0, 0, 0, 0, 0, 0, 0),
                (-97, 60, -96, 57, 64, -79, 19, 0, 0, 0, 0, 0, 0, 0, 0),
                (0, -170, 875, 231014, 643, 871, 89, 0, 0, 0, 0, 0, 0, 0, 0),
                (187, 64, 198, 64, 356087, 55, 484, 0, 0, 0, 0, 0, 0, 0, 0),
                (74, 174, 156, 63, 71, 576, 675, 0, 0, 0, 0, 0, 0, 0, 0),
                (362608, 362114, 363991, -475, 327, 432, 9, 0, 0, 0, 0, 0, 0, 0, 0),
                (193, 591, 1541, 889, 318875, 115, 130, 0, 0, 0, 0, 0, 0, 0, 0),
                (746, 602, 276, 552, 602, 576, 280, 0, 0, 0, 0, 0, 0, 0, 0),
                (38, 64, 180958, 64, 64, 704, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (64, 64, 170, 207, 429, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0)
                );
    constant children_left : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 13, 7, 9, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 13, 9, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1)
                );
    constant children_right : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 14, 8, 10, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 14, 10, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1)
                );
    constant value_int : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((0, 0, 0, 0, 0, 0, 0, 15, -72, -77, -107, 106, 74, 18, -80),
                (0, 0, 0, 0, 0, 0, 0, 49, -32, -71, -27, 66, -42, 4, -64),
                (0, 0, 0, 0, 0, 0, 0, 62, 39, 10, -43, -45, -66, 34, -29),
                (0, 0, 0, 0, 0, 0, 0, 29, -46, 51, -33, 51, 22, -1, -38),
                (0, 0, 0, 0, 0, 0, 0, 28, -43, -25, 14, -10, -44, -58, -33),
                (0, 0, 0, 0, 0, 0, 0, 9, -38, -16, -45, 32, -23, -11, -45),
                (0, 0, 0, 0, 0, 0, 0, 42, 21, -43, 26, 1, -26, 36, -18),
                (0, 0, 0, 0, 0, 0, 0, 11, -19, -42, -19, -38, -9, -52, -17),
                (0, 0, 0, 0, 0, 0, 0, 12, 33, 20, -4, -23, -50, 29, -11),
                (0, 0, 0, 0, 0, 0, 0, 13, -41, 13, -10, 46, 13, 24, -5),
                (0, 0, 0, 0, 0, 0, 0, -57, 1, -34, 10, 73, 1, -32, 17),
                (0, 0, 0, 0, 0, 0, 0, 4, -35, -55, -19, -27, -50, 32, -16),
                (0, 0, 0, 0, 0, 0, 0, 29, 4, -33, -2, 2, -18, 16, -9),
                (0, 0, 0, 0, 0, 0, 0, 27, -30, 8, -20, -11, -55, -43, 21),
                (0, 0, 0, 0, 0, 0, 0, 40, 15, -4, 5, -45, -20, 124, 0),
                (0, 0, 0, 0, 0, 0, 0, -31, 5, -21, 7, -33, -15, 3, -29),
                (0, 0, 0, 0, 0, 0, 0, 14, 53, 11, -2, 3, -5, 63, -17),
                (0, 0, 0, 0, 0, 0, 0, 3, -34, -33, 46, -74, -37, -3, -21),
                (0, 0, 0, 0, 0, 0, 0, 26, -12, 0, -77, 12, 40, -3, 4),
                (0, 0, 0, 0, 0, 0, 0, 9, -4, 0, 64, -49, -17, -20, 3),
                (0, 0, 0, 0, 0, 0, 0, -1, 18, -36, -1, -25, -93, -4, -38),
                (0, 0, 0, 0, 0, 0, 0, -27, -4, -13, 4, 3, 30, -33, 4),
                (0, 0, 0, 0, 0, 0, 0, -25, 5, 34, 4, -2, -44, 8, -5),
                (0, 0, 0, 0, 0, 0, 0, 1, -5, -21, 0, 44, -23, -21, 42),
                (0, 0, 0, 0, 0, 0, 0, 16, 51, 10, -5, 29, -7, -11, 6),
                (0, 0, 0, 0, 0, 0, 0, -52, 50, -82, -49, 4, -1, -24, 9),
                (0, 0, 0, 0, 0, 0, 0, -16, 2, 8, -1, -9, -38, -57, 2),
                (0, 0, 0, 0, 0, 0, 0, -16, 18, 6, -12, 3, -52, 19, -7),
                (0, 0, 0, 0, 0, 0, 0, 22, 4, 0, -18, -33, -16, 13, -29),
                (0, 0, 0, 0, 0, 0, 0, 34, -27, -10, 3, 12, -39, 4, -16),
                (0, 0, 0, 0, 0, 0, 0, 18, 0, -8, 2, 15, 36, -6, 29),
                (0, 0, 0, 0, 0, 0, 0, -34, 35, -3, 2, -56, -22, 0, -14),
                (0, 0, 0, 0, 0, 0, 0, 17, 56, -6, 10, 4, -1, -10, 0),
                (0, 0, 0, 0, 0, 0, 0, -33, 28, 34, 10, 0, -28, 6, -1),
                (0, 0, 0, 0, 0, 0, 0, -45, -8, 10, -1, 22, -25, -16, 2),
                (0, 0, 0, 0, 0, 0, 0, 7, -54, 0, 62, -48, 0, -2, -41),
                (0, 0, 0, 0, 0, 0, 0, -2, 9, -5, 2, 20, -33, -44, -16),
                (0, 0, 0, 0, 0, 0, 0, -13, 9, 17, 0, 0, 31, -10, 3),
                (0, 0, 0, 0, 0, 0, 0, -1, 3, 4, -34, 26, 68, 13, -35),
                (0, 0, 0, 0, 0, 0, 0, 11, 2, 0, -39, -50, 39, -2, 1),
                (0, 0, 0, 0, 0, 0, 0, -12, 2, 2, 22, 2, -3, 20, -18),
                (0, 0, 0, 0, 0, 0, 0, -22, 14, -16, 44, 0, 7, -4, 1),
                (0, 0, 0, 0, 0, 0, 0, 0, 13, -23, -4, -2, -19, 25, -25),
                (0, 0, 0, 0, 0, 0, 0, 40, -21, -12, 32, -1, 3, -14, 2),
                (0, 0, 0, 3, 0, 0, 0, -8, -63, 2, -1, -1, -16, 3, 3),
                (0, 0, 0, 0, 0, 0, 0, -3, 40, 3, -6, -15, 10, 1, -8),
                (0, 0, 0, 0, 0, 0, 0, -13, 1, -4, 3, 32, 6, -9, 1),
                (0, 0, 0, 0, 0, 0, 0, -12, 4, 44, -9, -32, 10, 1, -3),
                (0, 0, 0, 0, 0, 0, 0, -7, 3, 2, -17, 13, -8, 11, 4),
                (0, 0, 0, 0, 0, 0, 0, -14, 41, -54, 0, 0, 90, -52, -10),
                (0, 0, 0, 0, 0, 0, 0, -17, 21, 2, -4, -15, -65, 4, -4),
                (0, 0, 0, 0, 0, 0, 0, 4, -14, -1, -28, -9, 0, -2, 5),
                (0, 0, 0, 0, 0, 0, 0, 3, -17, 8, -2, 30, -6, -14, -47),
                (0, 0, 0, 0, 0, 0, 0, -23, 11, 6, -4, 2, -7, 20, 4),
                (0, 0, 0, 0, 0, 0, 0, 0, 3, 22, -22, -3, -27, 180, 13),
                (0, 0, 0, 0, 0, 0, 0, -36, -2, 0, -18, 15, -9, 14, -2),
                (0, 0, 0, 0, 0, 0, 0, 0, 31, -11, 38, 189, 25, -49, 13),
                (0, 0, 0, 0, 0, 0, 0, -42, 34, -50, 0, -4, 0, 12, -45),
                (0, 0, 0, 0, 0, 0, 0, -17, 23, -17, 2, -2, 3, 8, -10),
                (0, 0, 0, 0, 0, 0, 0, 16, 1, 2, -2, 6, -12, -11, -2),
                (0, 0, 0, 0, 0, 0, 0, -19, 0, 8, -1, 9, -13, -3, 13),
                (0, 0, 0, 0, 0, 0, 0, -6, 0, 20, 0, 24, -43, 0, -16),
                (0, 0, 0, 0, 0, 0, 0, -23, 13, -55, 34, -209, -14, -1, 1),
                (0, 0, 0, 0, 0, 0, 0, -8, 0, 16, 0, -6, 6, -1, -13),
                (0, 0, 0, 0, 0, 0, 0, -20, 18, 33, -32, 5, -26, 0, 3),
                (0, 0, 0, 0, 0, 0, 0, 11, -14, -18, 4, 11, -2, 1, -3),
                (0, 0, 0, 0, 0, 0, 0, 37, -23, -45, 11, -1, 1, -7, 77),
                (0, 0, 0, 0, 0, 0, 0, 17, -73, -1, 50, 0, -7, 3, -11),
                (0, 0, 0, 0, 0, 0, 0, -11, -58, 2, -19, 56, 5, -33, 0),
                (0, 0, 0, 0, 0, 0, 0, 23, -18, 61, 17, -4, 2, 3, 0),
                (0, 0, 0, 0, 0, 0, 0, 0, 51, 7, -9, -19, 6, 4, -11),
                (0, 0, 0, 0, 0, 0, 0, 0, -6, 3, -31, 0, -35, 11, -47),
                (0, 0, 0, 0, 0, 0, 0, -45, -9, 0, -8, -51, 28, 2, -25),
                (0, 0, 0, 0, 0, 0, 0, 11, 0, 2, -18, -1, -11, -4, 6),
                (0, 0, 0, 0, 0, 0, 0, -1, 1, -15, 6, 36, 5, -119, -3),
                (0, 0, 0, 0, 0, 0, 0, 22, -4, -32, 1, 3, -11, 1, -27),
                (0, 0, 0, 0, 93, 0, 0, -4, 0, -19, 14, -49, -11, 93, 93),
                (0, 0, 0, 0, 0, 0, 0, 47, 6, -5, 0, 13, -21, 59, -8),
                (0, 0, 0, 0, 0, 0, -32, 0, 36, -3, 10, 74, 0, -32, -32),
                (0, 0, 0, 0, 0, 0, 0, 0, 1, 1, -57, 117, 0, -24, 0),
                (0, 0, 0, 0, 0, 0, 0, -2, 2, 0, 7, 29, -34, -45, 0),
                (0, 0, 0, 0, 0, 0, 0, 0, -7, 4, -9, 19, 1, 1, -3),
                (0, 0, 0, 0, 0, 0, 0, -9, 3, -3, -17, 1, 10, 1, -26),
                (0, 0, 0, 0, 0, 0, 0, 0, -8, 25, -44, -23, 28, 3, -1),
                (0, 0, 0, 0, 0, 0, 0, -24, 13, -4, 0, -18, 2, 12, -1),
                (0, 0, 0, 0, 0, 0, 0, -2, 1, 0, 15, 13, -33, 142, 15),
                (0, 0, 0, 0, 0, 0, 0, 28, -44, 76, 15, 0, -127, 0, -5),
                (0, 0, 0, 0, 0, 0, 0, 38, 0, 11, 46, -5, -146, -9, 0),
                (0, 0, 0, 0, 0, 0, 0, -8, 33, -8, 2, 3, -14, -10, 0),
                (0, 0, 0, 0, 0, 0, 0, -3, 0, -40, 10, 14, -6, -9, 1),
                (0, 0, 0, 0, 0, 0, 0, -12, -135, 5, -8, -147, -13, -5, 0),
                (0, 0, 0, 0, 0, 0, 0, 0, -36, 12, -18, -125, -1, -5, 0),
                (0, 0, 0, 0, 0, 0, 0, 0, -99, 37, -21, 0, 38, 17, -18),
                (0, 0, 0, 0, 0, 0, 0, -26, 3, 19, -13, 5, -23, 1, -1),
                (0, 0, 0, 0, 0, 0, 0, -1, 10, 2, -18, 5, -5, -5, 4),
                (0, 0, 0, 0, 0, 0, 0, 31, 0, 15, -33, 2, 34, 29, 0),
                (0, 0, 0, 0, 0, 0, 0, 0, 4, 0, -10, -32, -2, 12, -36),
                (0, 0, 0, 0, 0, 0, 0, 0, 8, -71, -3, -5, 15, -40, -2),
                (0, 0, 0, 0, 0, 0, 0, 2, -2, 25, 1, -3, 4, -1, 5),
                (0, 0, 0, 0, 0, 0, 0, 11, 0, 7, -41, 5, -3, 12, 2)
                );
    constant parent : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 4, 4, 5, 5, 6, 6, 3, 3),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 5, 5, 6, 6, 4, 4),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6)
                );
    constant depth : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3)
                );
    constant iLeaf : intArray2D(nTrees-1 downto 0)(nLeaves-1 downto 0) := ((7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14)
                );
    constant value : tyArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := to_tyArray2D(value_int);
      constant threshold : txArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := to_txArray2D(threshold_int);
end Arrays0;