library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_misc.all;
  use ieee.numeric_std.all;

  use work.Constants.all;
  use work.Types.all;
  package Arrays0 is

    constant initPredict : ty := to_ty(0);
    constant feature : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((1, 0, 4, 4, 4, 19, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 4, 4, 3, 1, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 1, 0, 0, 17, 2, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 1, 0, 16, 3, 2, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 4, 4, 4, 16, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 3, 0, 17, 19, 0, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 1, 1, 4, 4, 4, 12, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 1, 1, 4, 4, 4, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 1, 1, 18, 4, 3, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 2, 4, 4, 17, 1, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 16, 0, 10, 18, 0, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 16, 18, 18, 1, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 20, 2, 13, 7, 16, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 18, 4, 4, 18, 1, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 1, 1, 2, 17, 5, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 16, 18, 18, 1, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 17, 2, 5, 16, 16, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 1, 18, 2, 0, 18, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 18, 4, 4, 0, 19, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 7, 3, 17, 6, 12, 14, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 2, 1, 6, 1, 17, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 17, 20, 7, 14, 16, 7, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 18, 16, 5, 16, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 4, 18, 19, 0, 3, 20, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 7, 12, 5, 6, 5, 15, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 16, 17, 17, 17, 7, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 20, 4, 10, 2, 1, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 3, 18, 4, 1, 16, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 7, 16, 12, 13, 10, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 17, 8, 7, 12, 17, 5, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 6, 17, 17, 2, 7, 12, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 1, 0, 5, 19, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 1, 4, 16, 16, 1, 20, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 16, 16, 20, 1, 2, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 6, 18, 17, 17, 16, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 18, 0, 19, 16, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 20, 14, 0, 5, 15, 13, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 4, 17, 5, 16, 17, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 17, 1, 19, 14, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 3, 16, 7, 20, 4, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 16, 2, 17, 2, 0, 5, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 18, 4, 20, 1, 18, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 17, 16, 5, 3, 3, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 4, 19, 6, 2, 10, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 2, 18, 4, 20, 18, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 16, 4, 2, 4, 20, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 1, 10, 19, 4, 6, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (7, 13, 13, 10, 12, 10, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 17, 17, 5, 17, 4, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 1, 16, 1, 16, 2, 19, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 0, 7, 4, 17, 13, 13, -2, -2, -2, -2, -2, -2, -2, -2),
                (6, 16, 17, 20, 2, 5, 10, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 17, 4, 18, 1, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 17, 8, 7, 14, 10, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 16, 0, 1, 6, 5, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 4, 3, 3, 3, 18, 19, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 17, 0, 8, 17, 4, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 6, 14, 20, 0, 12, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 7, 14, 5, 13, 15, 19, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 4, 17, 10, 10, 5, 10, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 4, 18, 2, 2, 4, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 0, 2, -2, -2, 5, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 17, 4, 20, 19, 0, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 19, 19, 16, 2, 14, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 6, 16, 0, 3, 2, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 13, 14, 5, 4, 15, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 9, 2, 10, 16, 4, 8, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 16, 2, 17, 5, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 16, 16, 8, 4, 16, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 18, 17, -2, 3, 20, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 19, 4, 13, 17, 10, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 2, 17, 0, 5, 16, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 2, 14, 12, 16, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (6, 16, 0, 4, 0, 3, 5, -2, -2, -2, -2, -2, -2, -2, -2),
                (19, 11, 17, 8, 1, 0, 12, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 4, 2, 3, 3, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 1, 10, 2, 15, 12, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 16, 3, 0, 20, 1, 7, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 16, 4, 4, 4, 1, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 7, 14, 5, 11, 15, 19, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 17, 9, 6, 2, 19, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 1, 4, 4, 2, 17, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 13, 13, 17, 4, 5, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (8, 10, 5, 16, 2, 7, 7, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 17, 17, 19, -2, 18, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 17, 9, 3, 2, 17, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 3, 17, 3, 0, 17, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 1, 18, 19, 17, -2, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 3, 0, 17, 19, 12, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 20, 6, 16, 11, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 8, 16, -2, 3, 4, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 3, 13, 18, 18, 3, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 12, 1, 3, 11, 19, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 17, 2, 16, 0, 18, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 1, 17, 5, 16, 1, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 20, 18, 19, 1, 5, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 1, 16, 16, -2, 6, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 18, 16, 0, 3, 2, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (5, 2, 2, 16, 17, 4, 9, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 4, 1, 4, 3, 0, -2, -2, -2, -2, -2, -2, -2, -2)
                );
    constant threshold_int : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((38848, 355904, 576, 576, 576, 320, 264128, 0, 0, 0, 0, 0, 0, 0, 0),
                (36928, 261952, 576, 576, 149184, 65984, 338240, 0, 0, 0, 0, 0, 0, 0, 0),
                (576, 24256, 386368, 317632, 52160, 261952, 457920, 0, 0, 0, 0, 0, 0, 0, 0),
                (576, 28992, 373056, 21952, 54080, 261952, 427072, 0, 0, 0, 0, 0, 0, 0, 0),
                (46272, 255424, 704, 576, 704, 34752, 364096, 0, 0, 0, 0, 0, 0, 0, 0),
                (576, 69184, 264384, 50752, 320, 169408, 155712, 0, 0, 0, 0, 0, 0, 0, 0),
                (211264, 73280, 26176, 576, 576, 704, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (190912, 50752, 58176, 576, 576, 704, 85312, 0, 0, 0, 0, 0, 0, 0, 0),
                (177216, 32064, 19520, 165568, 576, 135104, 50496, 0, 0, 0, 0, 0, 0, 0, 0),
                (112960, 261952, 704, 576, 57408, 15936, 193472, 0, 0, 0, 0, 0, 0, 0, 0),
                (576, 27072, 277440, 64, -145408, 118080, 111552, 0, 0, 0, 0, 0, 0, 0, 0),
                (68032, 120512, 38592, 181888, 157888, 97728, 54592, 0, 0, 0, 0, 0, 0, 0, 0),
                (704, 192, 261568, 64, 64, 23872, 473152, 0, 0, 0, 0, 0, 0, 0, 0),
                (84416, -147328, 704, 704, 139648, 13376, 177216, 0, 0, 0, 0, 0, 0, 0, 0),
                (93760, 29120, 15552, 24896, 15424, 64, 35648, 0, 0, 0, 0, 0, 0, 0, 0),
                (77120, 306752, 42944, -168448, -130048, 117184, -95488, 0, 0, 0, 0, 0, 0, 0, 0),
                (704, 14784, 261568, 64, 17728, 23488, 17088, 0, 0, 0, 0, 0, 0, 0, 0),
                (91584, 17472, 178048, 18112, 58560, -120448, 704, 0, 0, 0, 0, 0, 0, 0, 0),
                (103168, -93568, 576, 576, 292288, 320, 704, 0, 0, 0, 0, 0, 0, 0, 0),
                (71232, 64, 137280, 37568, 64, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (71616, 8896, 97856, 64, 25792, 49984, 45504, 0, 0, 0, 0, 0, 0, 0, 0),
                (78656, 70592, 576, 64, 64, 13120, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (13376, 169408, 162688, 23232, 64, 22976, 704, 0, 0, 0, 0, 0, 0, 0, 0),
                (-171328, 576, 93568, 320, 229888, 121536, 576, 0, 0, 0, 0, 0, 0, 0, 0),
                (49216, 64, 64, 64, 64, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (108736, 62912, 39488, 9920, 37824, 18368, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (47296, 576, 576, 64, 261952, 38336, 155392, 0, 0, 0, 0, 0, 0, 0, 0),
                (-197248, 249344, 198208, 704, 55360, 320, 371776, 0, 0, 0, 0, 0, 0, 0, 0),
                (122048, 64, 46912, 64, 64, 64, 200448, 0, 0, 0, 0, 0, 0, 0, 0),
                (57024, 33472, 64, 64, 64, 33600, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (101952, 64, 36160, 17600, 8896, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (260544, 8768, 387200, 64, 192, 46144, 30272, 0, 0, 0, 0, 0, 0, 0, 0),
                (47680, 117184, 576, 576, 34752, 30144, 704, 0, 0, 0, 0, 0, 0, 0, 0),
                (-212608, 46912, 14144, 192, 32448, 261952, 200128, 0, 0, 0, 0, 0, 0, 0, 0),
                (36416, 64, -72448, 80064, 24256, 46656, 80128, 0, 0, 0, 0, 0, 0, 0, 0),
                (260544, 211648, 384448, 192, 7744, 44608, 46144, 0, 0, 0, 0, 0, 0, 0, 0),
                (36160, 320, 64, 496192, 64, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (9408, 704, 23488, 64, 21696, 17344, 31424, 0, 0, 0, 0, 0, 0, 0, 0),
                (8128, 31424, 85696, 192, 64, 320, 38336, 0, 0, 0, 0, 0, 0, 0, 0),
                (5824, 132800, 12736, 64, 576, 704, 200128, 0, 0, 0, 0, 0, 0, 0, 0),
                (117184, 5824, 60096, 4416, 27968, 161728, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (47808, -212608, 576, 192, 126400, 127168, 17728, 0, 0, 0, 0, 0, 0, 0, 0),
                (4032, 23232, 46016, 64, 3392, 241216, 576, 0, 0, 0, 0, 0, 0, 0, 0),
                (11712, 576, 192, 64, 261952, 64, 33600, 0, 0, 0, 0, 0, 0, 0, 0),
                (576, 228800, 220288, 576, 704, -72448, 78656, 0, 0, 0, 0, 0, 0, 0, 0),
                (83968, 10816, 704, 261568, 576, 576, 364992, 0, 0, 0, 0, 0, 0, 0, 0),
                (126656, 38336, 64, 320, 576, 64, 27712, 0, 0, 0, 0, 0, 0, 0, 0),
                (64, 64, 64, 64, 64, 64, 704, 0, 0, 0, 0, 0, 0, 0, 0),
                (8768, 21952, 1344, 64, 37824, 704, 38336, 0, 0, 0, 0, 0, 0, 0, 0),
                (81984, 38336, 36288, 31424, 17600, 258624, 192, 0, 0, 0, 0, 0, 0, 0, 0),
                (320, 267328, 64, 576, 39424, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (64, 13760, 22592, 576, 149312, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (7488, 10432, 704, -106048, 34752, 14144, 27840, 0, 0, 0, 0, 0, 0, 0, 0),
                (59200, 31424, 64, 64, 64, 64, 23872, 0, 0, 0, 0, 0, 0, 0, 0),
                (73536, 36416, 32448, 8512, 38336, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (-171328, 576, 260544, 136128, 74816, 209728, 576, 0, 0, 0, 0, 0, 0, 0, 0),
                (47808, 9152, 104064, 64, 23744, 576, 156480, 0, 0, 0, 0, 0, 0, 0, 0),
                (71232, 64, 64, 576, 110528, 64, 55488, 0, 0, 0, 0, 0, 0, 0, 0),
                (39872, 64, 64, 64, 64, 64, 320, 0, 0, 0, 0, 0, 0, 0, 0),
                (13376, 576, 22464, 64, 64, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (-72448, 576, 80128, 128832, 256832, 576, 576, 0, 0, 0, 0, 0, 0, 0, 0),
                (192, 267328, 5824, 0, 0, 64, 142528, 0, 0, 0, 0, -256, -256, -256, -256),
                (47424, 87744, 576, 64, 448, 99136, 383744, 0, 0, 0, 0, 0, 0, 0, 0),
                (4032, 448, 320, 28608, 48832, 64, 30784, 0, 0, 0, 0, 0, 0, 0, 0),
                (-220288, 64, 832, 192576, 13376, 260992, 146624, 0, 0, 0, 0, 0, 0, 0, 0),
                (41536, 64, 64, 64, 704, 64, 43712, 0, 0, 0, 0, 0, 0, 0, 0),
                (90688, 64, 124480, 64, 29888, 704, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (140096, 3648, 139328, 1216, 64, 5568, 8768, 0, 0, 0, 0, 0, 0, 0, 0),
                (93504, 46016, 26880, 64, 576, 18752, 22976, 0, 0, 0, 0, 0, 0, 0, 0),
                (8512, -109376, 82496, 0, 832, 64, 49984, 0, 0, 0, 0, 0, 0, -256, -256),
                (38336, 320, 576, 64, 27712, 64, 704, 0, 0, 0, 0, 0, 0, 0, 0),
                (4928, 42176, 1344, 49856, 64, 9024, 38336, 0, 0, 0, 0, 0, 0, 0, 0),
                (117184, 5568, 64, 64, 832, 36288, 35520, 0, 0, 0, 0, 0, 0, 0, 0),
                (64, 26048, 313280, 576, 260160, 167744, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (192, 64, 30784, 64, 39232, 386496, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (32192, 576, 142528, 51904, 145600, 3904, 8768, 0, 0, 0, 0, 0, 0, 0, 0),
                (68032, 38336, 64, 25664, 64, 64, 704, 0, 0, 0, 0, 0, 0, 0, 0),
                (13248, 37824, 14656, 196032, 576, 38208, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (46016, 40896, 576, 576, 576, 28224, 178496, 0, 0, 0, 0, 0, 0, 0, 0),
                (42432, 64, 64, 64, 64, 64, 320, 0, 0, 0, 0, 0, 0, 0, 0),
                (23872, 17088, 64, 64, 17984, 192, 28608, 0, 0, 0, 0, 0, 0, 0, 0),
                (49984, 38336, 576, 576, 147264, 58560, 440448, 0, 0, 0, 0, 0, 0, 0, 0),
                (39360, 64, 64, 33600, 576, 64, 74176, 0, 0, 0, 0, 0, 0, 0, 0),
                (64, 64, 64, 26304, 261952, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (320, 38912, 94912, 192, 0, 80128, 31872, 0, 0, 0, 0, 0, 0, -256, -256),
                (23872, 17344, 64, 45632, 24128, 26304, 8256, 0, 0, 0, 0, 0, 0, 0, 0),
                (-212608, 153152, 82112, 76352, 386112, 79680, -54208, 0, 0, 0, 0, 0, 0, 0, 0),
                (93632, 2368, -148800, 320, 39360, 0, 151616, 0, 0, 0, 0, 0, 0, -256, -256),
                (47808, 260544, 336960, 22464, 576, 64, 255552, 0, 0, 0, 0, 0, 0, 0, 0),
                (126400, 8512, 192, 64, 704, 64, 32192, 0, 0, 0, 0, 0, 0, 0, 0),
                (192, 64, 4288, 0, 67328, 576, 201536, 0, 0, 0, 0, 0, 0, -256, -256),
                (220288, 2368, 64, -8128, -68608, 155648, 16128, 0, 0, 0, 0, 0, 0, 0, 0),
                (39360, 64, 21568, 212544, 64, 448, 20288, 0, 0, 0, 0, 0, 0, 0, 0),
                (82496, 79936, 34880, 46016, 178496, 57088, -53248, 0, 0, 0, 0, 0, 0, 0, 0),
                (1472, 43072, 1600, 64, 44416, 45376, 320, 0, 0, 0, 0, 0, 0, 0, 0),
                (-212608, 576, -211648, 320, 18176, 64, 94016, 0, 0, 0, 0, 0, 0, 0, 0),
                (155328, 153920, 40640, 47936, 0, 64, 311744, 0, 0, 0, 0, 0, 0, -256, -256),
                (56128, 18688, 4288, 409280, 260864, 261824, 72768, 0, 0, 0, 0, 0, 0, 0, 0),
                (64, 139712, 70080, 29888, 19904, 576, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (38336, 408640, 576, 32576, 704, 141248, 440448, 0, 0, 0, 0, 0, 0, 0, 0)
                );
    constant children_left : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 11, 13, 7, 9, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 13, 7, 9, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 13, 9, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 13, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 13, 7, 9, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 13, 9, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1)
                );
    constant children_right : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 12, 14, 8, 10, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 14, 8, 10, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 14, 10, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 14, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 14, 8, 10, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 14, 10, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1)
                );
    constant value_int : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((0, 0, 0, 0, 0, 0, 0, 24, 61, -37, 9, -57, -27, 60, -9),
                (0, 0, 0, 0, 0, 0, 0, 38, 52, 26, -27, -31, -49, 34, -27),
                (0, 0, 0, 0, 0, 0, 0, 26, -17, -36, 0, 44, 27, -2, -30),
                (0, 0, 0, 0, 0, 0, 0, -16, 21, -12, -36, 40, 22, 5, -21),
                (0, 0, 0, 0, 0, 0, 0, 25, 37, -1, 25, -33, -11, 27, -12),
                (0, 0, 0, 0, 0, 0, 0, -3, 34, -30, -5, 36, 29, 16, -17),
                (0, 0, 0, 0, 0, 0, 0, 21, 33, -27, 20, 4, 21, -25, -3),
                (0, 0, 0, 0, 0, 0, 0, 20, 31, -14, 24, -1, 17, -18, -33),
                (0, 0, 0, 0, 0, 0, 0, 28, -9, -5, 24, 14, -10, -14, 9),
                (0, 0, 0, 0, 0, 0, 0, 8, 27, -3, 25, -6, -24, 11, -20),
                (0, 0, 0, 0, 0, 0, 0, -13, -35, -34, 10, 28, 18, 9, -6),
                (0, 0, 0, 0, 0, 0, 0, 24, -28, 4, -32, -19, -33, 13, -13),
                (0, 0, 0, 0, 0, 0, 0, -19, 20, -23, 2, 31, 18, 9, -17),
                (0, 0, 0, 0, 0, 0, 0, -31, 16, 10, -20, -1, -17, 10, -12),
                (0, 0, 0, 0, 0, 0, 0, 27, 18, -9, 20, 17, 5, -10, 3),
                (0, 0, 0, 0, 0, 0, 0, -27, 9, -21, -2, -18, -32, -22, 14),
                (0, 0, 0, 0, 0, 0, 0, 14, -22, -9, 6, 28, 12, 10, 0),
                (0, 0, 0, 0, 0, 0, 0, 26, 19, 17, 1, -15, 2, -31, 11),
                (0, 0, 0, 0, 0, 0, 0, -15, 2, 9, 0, -23, -4, -5, 10),
                (0, 0, 0, 0, 0, 0, 0, -36, 2, -21, 7, -20, 21, 12, -6),
                (0, 0, 0, 0, 0, 0, 0, 8, 27, 16, 5, -2, 7, -24, 15),
                (0, 0, 0, 0, 0, 0, 0, -6, 6, 29, 11, -18, -6, -31, 6),
                (0, 0, 0, 0, 0, 0, 0, 23, 10, 12, 1, -6, 2, -22, 7),
                (0, 0, 0, 0, 0, 0, 0, -26, -6, 16, -9, 3, -5, -10, 8),
                (0, 0, 0, 0, 0, 0, 0, 20, -19, -16, 5, 4, -36, 20, 0),
                (0, 0, 0, 0, 0, 0, 0, 3, 17, -2, 4, -30, -20, -17, 14),
                (0, 0, 0, 0, 0, 0, 0, 0, -23, 11, 0, 20, 46, -6, 32),
                (0, 0, 0, 0, 0, 0, 0, -25, 15, 12, -22, -51, 1, -24, -4),
                (0, 0, 0, 0, 0, 0, 0, -21, 4, 5, -13, -20, -34, 49, 0),
                (0, 0, 0, 0, 0, 0, 0, -24, 3, -10, 10, -14, -2, 17, -1),
                (0, 0, 0, 0, 0, 0, 0, -25, 5, 22, 7, -19, 0, -14, 4),
                (0, 0, 0, 0, 0, 0, 0, 13, 4, 2, -2, -29, 6, -12, 5),
                (0, 0, 0, 0, 0, 0, 0, -32, 0, -23, -7, 20, 39, 3, -48),
                (0, 0, 0, 0, 0, 0, 0, -8, -25, 0, 46, 14, -8, -3, 3),
                (0, 0, 0, 0, 0, 0, 0, -8, 24, 23, 9, -4, 9, 2, -4),
                (0, 0, 0, 0, 0, 0, 0, 3, -1, 7, -23, -25, -1, -5, 24),
                (0, 0, 0, 0, 0, 0, 0, -16, 80, 12, -1, 14, -10, -17, 2),
                (0, 0, 0, 0, 0, 0, 0, 6, -13, 14, -5, 1, 12, -7, 1),
                (0, 0, 0, 0, 0, 0, 0, 4, -18, 23, 2, -41, 0, -15, 6),
                (0, 0, 0, 0, 0, 0, 0, 7, 21, -24, 17, -9, 8, -3, 2),
                (0, 0, 0, 0, 0, 0, 0, 0, 28, 8, -1, 1, -21, 3, -1),
                (0, 0, 0, 0, 0, 0, 0, -2, -20, 0, -15, 25, -7, 12, -16),
                (0, 0, 0, 0, 0, 0, 0, 28, 10, 24, 1, 0, -6, 14, -5),
                (0, 0, 0, 0, 0, 0, 0, -24, -3, 9, -2, 9, -4, -8, 1),
                (0, 0, 0, 0, 0, 0, 0, -20, 32, -37, 0, -2, 1, -19, 33),
                (0, 0, 0, 0, 0, 0, 0, 13, -7, 4, -1, -6, 3, 8, -11),
                (0, 0, 0, 0, 0, 0, 0, -2, 2, 6, -4, -21, -4, -9, -33),
                (0, 0, 0, 0, 0, 0, 0, -18, 8, -12, 5, 6, -2, -21, 2),
                (0, 0, 0, 0, 0, 0, 0, 21, 4, -3, 3, -13, 2, -1, 2),
                (0, 0, 0, 0, 0, 0, 0, 0, -5, -5, 5, -18, -7, 15, -6),
                (0, 0, 0, 0, 0, 0, 0, -17, 22, -28, -54, -9, 2, 2, -5),
                (0, 0, 0, 0, 0, 0, 0, -17, 7, -10, 3, 10, 1, 0, -16),
                (0, 0, 0, 0, 0, 0, 0, -38, -5, 3, 15, -5, 0, 6, -4),
                (0, 0, 0, 0, 0, 0, 0, -10, 0, 7, 1, -2, -21, 3, -6),
                (0, 0, 0, 0, 0, 0, 0, 29, 8, 0, 2, -16, -5, -9, 6),
                (0, 0, 0, 0, 0, 0, 0, -13, 3, 9, -4, 1, -12, -2, -19),
                (0, 0, 0, 0, 0, 0, 0, -16, -1, 3, 0, 29, 7, 3, 27),
                (0, 0, 0, 0, 0, 0, 0, -7, 12, 4, 0, -32, 14, 12, -1),
                (0, 0, 0, 0, 0, 0, 0, 28, -13, 1, -5, 15, -10, -15, 1),
                (0, 0, 0, 0, 0, 0, 0, -1, -16, -12, 3, 17, 2, 0, -10),
                (0, 0, 0, 0, 0, 0, 0, -10, -2, 6, -2, 3, 0, -4, 1),
                (0, 0, 0, -5, -36, 0, 0, -5, 12, -2, 0, -5, -5, -36, -36),
                (0, 0, 0, 0, 0, 0, 0, -5, 0, 50, 8, 24, 7, -5, 21),
                (0, 0, 0, 0, 0, 0, 0, 10, 1, 18, -8, 0, -12, 3, -4),
                (0, 0, 0, 0, 0, 0, 0, -31, 20, 6, -20, 23, -27, 0, -14),
                (0, 0, 0, 0, 0, 0, 0, 6, -1, -14, 4, 14, -8, 13, -2),
                (0, 0, 0, 0, 0, 0, 0, 2, -14, 2, -6, -12, 4, -2, 3),
                (0, 0, 0, 0, 0, 0, 0, -13, 27, -8, 3, 21, -7, -3, 1),
                (0, 0, 0, 0, 0, 0, 0, -1, 1, 9, -3, 25, -21, 3, 39),
                (0, 0, 0, -2, 0, 0, 0, 8, 35, -5, 0, 6, -9, -2, -2),
                (0, 0, 0, 0, 0, 0, 0, -1, -7, -11, 2, 7, -14, -8, 3),
                (0, 0, 0, 0, 0, 0, 0, -3, 18, 8, 1, -15, -2, 0, 1),
                (0, 0, 0, 0, 0, 0, 0, 12, -5, -9, 0, -20, -2, 27, -7),
                (0, 0, 0, 0, 0, 0, 0, -11, 1, -6, 4, 1, -15, 3, -2),
                (0, 0, 0, 0, 0, 0, 0, -7, 1, 10, 35, -7, 17, -5, 1),
                (0, 0, 0, 0, 0, 0, 0, 2, -12, 11, -12, 22, -3, -2, 1),
                (0, 0, 0, 0, 0, 0, 0, 5, 0, 4, -7, 4, -4, -15, 4),
                (0, 0, 0, 0, 0, 0, 0, 9, 1, 1, -10, -1, 7, -2, 0),
                (0, 0, 0, 0, 0, 0, 0, -1, 1, 2, -5, 3, 13, -4, 14),
                (0, 0, 0, 0, 0, 0, 0, 22, -8, -1, 3, 13, -5, -8, 1),
                (0, 0, 0, 0, 0, 0, 0, -7, 1, 19, 4, 6, -1, -17, -5),
                (0, 0, 0, 0, 0, 0, 0, -1, 1, -5, 5, 2, -9, -9, 11),
                (0, 0, 0, 0, 0, 0, 0, 0, 8, -18, -1, -20, 3, 3, -1),
                (0, 0, 0, 0, 0, 0, 0, -2, 1, -2, -24, 47, 0, -7, 1),
                (0, 0, 0, 0, -39, 0, 0, -15, 12, 0, -1, 7, 39, -39, -39),
                (0, 0, 0, 0, 0, 0, 0, -3, 1, 16, 3, 9, 0, 5, -7),
                (0, 0, 0, 0, 0, 0, 0, -6, -24, 36, -2, 0, -9, -4, 6),
                (0, 0, 0, 0, 0, 37, 0, 9, -5, 0, 1, -9, 32, 37, 37),
                (0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -16, 16, 3, 28, -16),
                (0, 0, 0, 0, 0, 0, 0, -2, 30, -9, 0, 36, -11, 5, -16),
                (0, 0, 0, -32, 0, 0, 0, 1, -23, -15, 9, -2, 0, -32, -32),
                (0, 0, 0, 0, 0, 0, 0, 10, -2, -1, 0, -23, 15, 40, 0),
                (0, 0, 0, 0, 0, 0, 0, 1, -5, -11, -1, 4, 0, 5, -2),
                (0, 0, 0, 0, 0, 0, 0, 0, 2, 12, -8, 22, -1, -5, 4),
                (0, 0, 0, 0, 0, 0, 0, 9, -2, -14, 17, 23, -15, -18, 0),
                (0, 0, 0, 0, 0, 0, 0, -15, 3, 39, 0, -4, 50, 0, 19),
                (0, 0, 0, 0, 34, 0, 0, 0, 8, -30, -9, 19, -14, 34, 34),
                (0, 0, 0, 0, 0, 0, 0, 0, 3, 2, -7, 27, 0, -1, -6),
                (0, 0, 0, 0, 0, 0, 0, -23, -1, 11, 1, -2, 6, 0, -3),
                (0, 0, 0, 0, 0, 0, 0, 0, -4, 7, -6, 5, -7, -4, 9)
                );
    constant parent : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 5, 5, 6, 6, 3, 3, 4, 4),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 4, 4, 5, 5, 6, 6, 3, 3),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 5, 5, 6, 6, 4, 4),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 6, 6, 5, 5),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 4, 4, 5, 5, 6, 6, 3, 3),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 5, 5, 6, 6, 4, 4),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6)
                );
    constant depth : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3)
                );
    constant iLeaf : intArray2D(nTrees-1 downto 0)(nLeaves-1 downto 0) := ((7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14)
                );
    constant value : tyArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := to_tyArray2D(value_int);
      constant threshold : txArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := to_txArray2D(threshold_int);
end Arrays0;