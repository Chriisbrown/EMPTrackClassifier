library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_misc.all;
  use ieee.numeric_std.all;

  use work.Constants.all;
  use work.Types.all;
  package Arrays0 is

    constant initPredict : ty := to_ty(0);
    constant feature : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((4, 1, 0, 3, 1, 0, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 1, 0, 0, 19, 3, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 4, 4, 3, 1, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 17, 0, 0, 3, 0, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 1, 3, 0, 3, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 3, 4, 0, 4, 18, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 17, 5, 4, 4, 12, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 1, 4, 17, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 3, 4, 0, 16, 18, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 7, 17, 17, 6, 16, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 17, 1, 7, 13, 3, 20, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 0, 20, 18, 20, 15, 7, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 3, 18, 17, 16, 1, 20, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 1, 16, 5, 16, 9, 12, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 2, 4, 6, 5, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 17, 4, 7, 19, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 1, 2, 5, 17, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 0, 1, 20, 16, 18, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 7, 4, 12, 13, 1, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 4, 4, 16, 16, 16, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 0, 0, 4, 1, 16, 20, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 17, 8, 20, 14, 10, 5, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 2, 16, 4, 17, 14, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (7, 13, 6, 10, 12, 20, 13, -2, -2, -2, -2, -2, -2, -2, -2),
                (10, 17, 4, 5, 19, 7, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 1, 15, 16, 5, 17, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (14, 17, 19, 7, 15, 0, 13, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 16, 17, 16, 4, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 2, 3, 4, 3, 1, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (6, 16, 0, 4, 0, 16, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 5, 10, 7, 2, 3, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 4, 1, 16, 16, 17, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 0, 3, 17, 7, 12, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 4, 3, 0, 3, 3, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 1, 1, 17, 19, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 1, 17, 3, 3, 16, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 20, 14, 20, 17, 16, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 3, 17, 18, 17, 4, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 5, 16, 17, 16, 17, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 4, 1, 17, 16, 3, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 13, 10, 3, 2, 20, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 17, 9, 2, 4, 19, 6, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 1, 1, 2, 1, 1, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 1, 16, 16, 20, 4, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 2, 0, 16, 16, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 4, 0, 3, 0, 16, 5, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 2, 16, 16, 16, 2, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 20, 12, 11, 12, 5, 19, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 0, 20, 4, 17, 2, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 17, 4, 17, 17, 0, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 16, 3, 20, 2, 2, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 12, 1, 6, 14, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (20, 4, 5, 12, 2, 2, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 16, 16, 16, 14, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 4, 19, 16, 16, 13, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 20, 0, 16, 17, 1, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 20, 3, 1, 3, 9, 20, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 17, 16, 18, 0, -2, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 4, 18, 14, 3, 4, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 7, 17, 5, 13, 3, 13, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 16, 2, 3, 1, 3, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 16, 1, 16, -2, 16, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 17, 1, 3, -2, 0, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (10, 20, 2, 17, 16, 4, 8, -2, -2, -2, -2, -2, -2, -2, -2),
                (11, 7, 7, 5, 17, 17, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 20, 12, 6, 3, 4, 15, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 19, 19, 6, 0, 6, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 16, 2, 4, 0, 14, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (20, 2, 17, 16, 16, 0, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 2, 0, 4, 4, 4, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 4, 1, 2, 2, 2, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (8, 2, 3, 17, 10, 6, 6, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 0, 3, 0, 1, 16, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 20, 1, 18, 0, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 16, 1, 18, 6, 10, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 2, 17, 4, 5, 2, 20, -2, -2, -2, -2, -2, -2, -2, -2),
                (14, 17, 2, 15, 0, 17, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 3, 0, 18, 4, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 3, 3, 17, 8, 18, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 16, 17, 3, 3, 6, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 2, 16, 17, 16, 2, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 16, 16, 4, 4, 17, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 2, 16, 17, 17, 18, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 3, 3, 3, 18, 3, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 16, 16, 1, 3, 3, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 1, 1, 0, 17, 16, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 0, 0, 4, 0, 4, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 0, 0, 16, 16, 4, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (20, 19, 0, 2, 17, 3, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 3, 2, 0, 1, 4, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 1, 3, 10, 10, 16, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 0, 1, 2, 3, 18, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 17, 0, 17, 15, 13, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 3, 14, 3, 2, 18, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 14, 0, 6, 16, 18, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 16, 18, 1, 17, 1, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 17, 2, 16, 18, 17, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 16, 16, 1, 2, 3, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 1, 0, 3, 5, 16, 20, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 17, 1, 18, 2, 16, 0, -2, -2, -2, -2, -2, -2, -2, -2)
                );
    constant threshold_int : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((576, 53, 426, 178, 115, 348, 260, 0, 0, 0, 0, 0, 0, 0, 0),
                (576, 73, 487, 304, 320, 292, 71, 0, 0, 0, 0, 0, 0, 0, 0),
                (106, 379, 704, 576, 233, 161, 368, 0, 0, 0, 0, 0, 0, 0, 0),
                (576, 412, 319, 210, 204, 256, 704, 0, 0, 0, 0, 0, 0, 0, 0),
                (126, 581, 188, 267, 730, 192, 302212, 0, 0, 0, 0, 0, 0, 0, 0),
                (1061, 226, 704, 260, 704, 1264, 308, 0, 0, 0, 0, 0, 0, 0, 0),
                (18, 634, 453, 64, 576, 704, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (165, 281, 218, 576, 388, 254329, 293518, 0, 0, 0, 0, 0, 0, 0, 0),
                (941, 296, 576, 763, 248994, 1376, 231, 0, 0, 0, 0, 0, 0, 0, 0),
                (200, 64, 134, 290, 64, 308205, 233, 0, 0, 0, 0, 0, 0, 0, 0),
                (191, 549, -3, 64, 64, 333, 704, 0, 0, 0, 0, 0, 0, 0, 0),
                (55, 261, 192, 1586, 576, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (1331, 329, 1639, 277, 217314, -40, 576, 0, 0, 0, 0, 0, 0, 0, 0),
                (678, 228, 20681, 64, 305900, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (694, -2, 704, 64, 64, 162879, 213363, 0, 0, 0, 0, 0, 0, 0, 0),
                (137, 110, 704, 64, 192, 162154, 174635, 0, 0, 0, 0, 0, 0, 0, 0),
                (811, -85, 844, 64, 92, 20681, 16960, 0, 0, 0, 0, 0, 0, 0, 0),
                (-71, 323, 253, 576, 363234, 1534, 264242, 0, 0, 0, 0, 0, 0, 0, 0),
                (373673, 64, 576, 64, 64, 50, 164, 0, 0, 0, 0, 0, 0, 0, 0),
                (453, 704, 704, 134920, 223571, 217347, 564, 0, 0, 0, 0, 0, 0, 0, 0),
                (4248, 404, 834, 576, 59, 21340, 704, 0, 0, 0, 0, 0, 0, 0, 0),
                (42, 249, 64, 320, 64, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (264, 98, 343409, 576, 276, 64, 42, 0, 0, 0, 0, 0, 0, 0, 0),
                (64, 64, 64, 64, 64, 576, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (64, 86, 576, 64, 192, 64, 127840, 0, 0, 0, 0, 0, 0, 0, 0),
                (-157, 147, 64, 140518, 64, 376, 576, 0, 0, 0, 0, 0, 0, 0, 0),
                (64, 332, 320, 64, 64, 152, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (789, 371434, 141, 308304, 576, 57663, 29013, 0, 0, 0, 0, 0, 0, 0, 0),
                (5071, 369, 434, 576, 450, 74, 704, 0, 0, 0, 0, 0, 0, 0, 0),
                (64, 176018, 350, 576, 390, 53415, 246, 0, 0, 0, 0, 0, 0, 0, 0),
                (185, 64, 64, 64, 295, 159, 138, 0, 0, 0, 0, 0, 0, 0, 0),
                (566, 576, -35, 161035, 230849, 178, 361291, 0, 0, 0, 0, 0, 0, 0, 0),
                (1721, -51, 444, 41, 64, 64, 88, 0, 0, 0, 0, 0, 0, 0, 0),
                (844, 704, 201, 486, 318, 194, 144437, 0, 0, 0, 0, 0, 0, 0, 0),
                (-155, 59, -139, 245, 320, 182341, 6981, 0, 0, 0, 0, 0, 0, 0, 0),
                (275, 72, 263, 231, 89, 16103, 145, 0, 0, 0, 0, 0, 0, 0, 0),
                (275, 320, 64, 192, 134, 103964, 576, 0, 0, 0, 0, 0, 0, 0, 0),
                (374562, 468, 640, 1751, 558, 704, -4, 0, 0, 0, 0, 0, 0, 0, 0),
                (211, 64, 254757, 170, 278929, 141, 409, 0, 0, 0, 0, 0, 0, 0, 0),
                (14, 576, 106, 126, 307283, 260, 258116, 0, 0, 0, 0, 0, 0, 0, 0),
                (-206, 64, 64, 423, 138, 576, 576, 0, 0, 0, 0, 0, 0, 0, 0),
                (179, 136, 64, 524, 704, 192, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (2503, 59, 146, 365, 81, 119, 504, 0, 0, 0, 0, 0, 0, 0, 0),
                (-216, 147, 147961, 122637, 576, 576, 576, 0, 0, 0, 0, 0, 0, 0, 0),
                (704, 313, 637, 31614, 23546, 84436, 59309, 0, 0, 0, 0, 0, 0, 0, 0),
                (89, 704, 264, 248, 128, 74787, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (187, 436, 198774, 34413, 228643, 647, 424, 0, 0, 0, 0, 0, 0, 0, 0),
                (299, 320, 64, 64, 64, 64, 320, 0, 0, 0, 0, 0, 0, 0, 0),
                (78311, 409, 576, 576, 421, 477, 254823, 0, 0, 0, 0, 0, 0, 0, 0),
                (362970, 186, 576, 134, 220, 681, 294, 0, 0, 0, 0, 0, 0, 0, 0),
                (704, 59079, 313, 576, 473, 158, 593, 0, 0, 0, 0, 0, 0, 0, 0),
                (103, 64, -34, 64, 64, 308666, 257787, 0, 0, 0, 0, 0, 0, 0, 0),
                (64, 576, 64, 64, 475, 171, 72, 0, 0, 0, 0, 0, 0, 0, 0),
                (253, 329, 264242, 34282, 10769, 64, 214, 0, 0, 0, 0, 0, 0, 0, 0),
                (574, 576, 320, 259862, 279061, 64, 96, 0, 0, 0, 0, 0, 0, 0, 0),
                (638, 64, 668, 84601, 625, 42, 172001, 0, 0, 0, 0, 0, 0, 0, 0),
                (97, 704, 260, 194, -73, 64, 576, 0, 0, 0, 0, 0, 0, 0, 0),
                (306, 2, 55292, 139, -89, 0, 344, 0, 0, 0, 0, 0, 0, -256, -256),
                (101, 576, 139, 64, 100, 576, 704, 0, 0, 0, 0, 0, 0, 0, 0),
                (296, 64, 421, 64, 64, 196, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (369425, 369030, 515, 477, 42, 361, 576, 0, 0, 0, 0, 0, 0, 0, 0),
                (-598, 369128, -313, 229236, 0, 83086, -289, 0, 0, 0, 0, 0, 0, -256, -256),
                (2503, 560, -170, -88, 0, 801, -168, 0, 0, 0, 0, 0, 0, -256, -256),
                (64, 576, 548, 200, 200157, 576, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (64, 64, 64, 64, 208, 293, 576, 0, 0, 0, 0, 0, 0, 0, 0),
                (245, 320, 64, 64, 173, 576, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (359, 576, 576, 64, 495, 64, 685, 0, 0, 0, 0, 0, 0, 0, 0),
                (639, 245010, 220, 576, 691, 64, 212045, 0, 0, 0, 0, 0, 0, 0, 0),
                (704, 577, 81, 245142, 17651, 545, 789, 0, 0, 0, 0, 0, 0, 0, 0),
                (18507, 420, 424, 576, 576, 576, 415, 0, 0, 0, 0, 0, 0, 0, 0),
                (15478, 576, 20, 730, 505, 638, 125, 0, 0, 0, 0, 0, 0, 0, 0),
                (64, 135, 188, 179, 64, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (811, 807, 201, 807, 165, 154811, 559, 0, 0, 0, 0, 0, 0, 0, 0),
                (264, 859, 192, -243, 836, 601, 314232, 0, 0, 0, 0, 0, 0, 0, 0),
                (-312, 275373, -34, 229, 64, 64, 20, 0, 0, 0, 0, 0, 0, 0, 0),
                (94, 168, 95, 576, 64, 241, 704, 0, 0, 0, 0, 0, 0, 0, 0),
                (64, 558, 163, 64, 803, 456, 576, 0, 0, 0, 0, 0, 0, 0, 0),
                (341, 340, 432, 1766, 704, 274944, 224757, 0, 0, 0, 0, 0, 0, 0, 0),
                (505, 208, 201, 330, 64, 1121, 306, 0, 0, 0, 0, 0, 0, 0, 0),
                (17, 41000, 19, 244, 286, 64, 106, 0, 0, 0, 0, 0, 0, 0, 0),
                (7179, 563, 13831, 150, 3886, 400, 14226, 0, 0, 0, 0, 0, 0, 0, 0),
                (487, 40901, 94480, 576, 576, 517, 303035, 0, 0, 0, 0, 0, 0, 0, 0),
                (35500, 403, 36554, 133, 54, 836, 83, 0, 0, 0, 0, 0, 0, 0, 0),
                (568, 455, 177, 401, 1549, -56, 874, 0, 0, 0, 0, 0, 0, 0, 0),
                (362970, 362773, 363793, 147, 58, 235, 576, 0, 0, 0, 0, 0, 0, 0, 0),
                (-384, -500, -370, 362, 236, 217940, 704, 0, 0, 0, 0, 0, 0, 0, 0),
                (1024, 205, 231, 576, 232, 576, 789, 0, 0, 0, 0, 0, 0, 0, 0),
                (174, 171, 211, 18244, 212375, 576, 218, 0, 0, 0, 0, 0, 0, 0, 0),
                (704, 192, 629, 582, 223, 109, 193, 0, 0, 0, 0, 0, 0, 0, 0),
                (266283, 158, 689, 607, 33, 576, 230, 0, 0, 0, 0, 0, 0, 0, 0),
                (704, 57, 39, 64, 64, 112099, 650, 0, 0, 0, 0, 0, 0, 0, 0),
                (740, 740, 126, 738, -30, 1309, 322, 0, 0, 0, 0, 0, 0, 0, 0),
                (566, 715, 604, 700, 64, 64, 336658, 0, 0, 0, 0, 0, 0, 0, 0),
                (575, 549, 64, 548, 278, 671, -41, 0, 0, 0, 0, 0, 0, 0, 0),
                (179, 64, 181, 64, 154679, 161, 374924, 0, 0, 0, 0, 0, 0, 0, 0),
                (375056, 374924, 56, 106, 52, -131, 377, 0, 0, 0, 0, 0, 0, 0, 0),
                (-230, 173, -228, 152242, 514, 134, -65, 0, 0, 0, 0, 0, 0, 0, 0),
                (71, 176348, 197819, 31, 493, 196, 380, 0, 0, 0, 0, 0, 0, 0, 0),
                (196, 106, 490, 172, 64, 70276, 320, 0, 0, 0, 0, 0, 0, 0, 0),
                (48936, 496, 143, 641, 554, 49430, 382, 0, 0, 0, 0, 0, 0, 0, 0)
                );
    constant children_left : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 13, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 13, 9, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 13, 9, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1)
                );
    constant children_right : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 14, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 14, 10, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 14, 10, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1)
                );
    constant value_int : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((0, 0, 0, 0, 0, 0, 0, 15, -73, -74, -107, 105, 71, 19, -80),
                (0, 0, 0, 0, 0, 0, 0, 58, -34, -73, -36, 66, -42, 5, -56),
                (0, 0, 0, 0, 0, 0, 0, 27, 57, 7, -44, -42, -66, 51, -12),
                (0, 0, 0, 0, 0, 0, 0, 29, -45, 60, -30, 55, 40, -16, 24),
                (0, 0, 0, 0, 0, 0, 0, 29, -25, -11, -42, -12, -47, -58, -36),
                (0, 0, 0, 0, 0, 0, 0, 37, 8, -34, 4, -36, -59, 24, -48),
                (0, 0, 0, 0, 0, 0, 0, 44, 15, -28, 0, -29, 9, -47, 29),
                (0, 0, 0, 0, 0, 0, 0, 7, 33, -8, 18, -33, -3, -54, -25),
                (0, 0, 0, 0, 0, 0, 0, 11, -26, -39, -13, -31, -52, 42, -8),
                (0, 0, 0, 0, 0, 0, 0, -61, 7, -39, 14, -51, -15, -8, -36),
                (0, 0, 0, 0, 0, 0, 0, -9, 10, -31, 35, 6, -25, -22, 2),
                (0, 0, 0, 0, 0, 0, 0, 31, -38, -24, 34, 36, -4, -17, -1),
                (0, 0, 0, 0, 0, 0, 0, -2, 11, -33, -7, 3, -27, -45, -18),
                (0, 0, 0, 0, 0, 0, 0, 15, 0, -42, 2, -70, -44, -21, -3),
                (0, 0, 0, 0, 0, 0, 0, 9, 31, 13, 0, -26, -7, 21, -12),
                (0, 0, 0, 0, 0, 0, 0, -44, -5, 21, 6, -22, -4, 22, -9),
                (0, 0, 0, 0, 0, 0, 0, 27, 6, -9, 1, -62, -16, -73, -36),
                (0, 0, 0, 0, 0, 0, 0, 18, 38, -40, 26, 0, -24, -48, -12),
                (0, 0, 0, 0, 0, 0, 0, -37, 5, 7, -20, 48, 104, -39, 15),
                (0, 0, 0, 0, 0, 0, 0, -14, 3, 16, -11, -31, 3, -4, -55),
                (0, 0, 0, 0, 0, 0, 0, -56, 56, -88, -45, 16, 0, -18, -44),
                (0, 0, 0, 0, 0, 0, 0, -34, 1, 31, 1, -3, -47, 36, -2),
                (0, 0, 0, 0, 0, 0, 0, -4, 19, -3, 3, -46, -17, 91, -20),
                (0, 0, 0, 0, 0, 0, 0, -36, 3, -29, 10, -29, 18, 8, -11),
                (0, 0, 0, 0, 0, 0, 0, 22, -21, 17, -1, 12, -52, 18, -11),
                (0, 0, 0, 0, 0, 0, 0, -5, 33, -53, 13, -2, 15, -34, 0),
                (0, 0, 0, 0, 0, 0, 0, -17, 2, 40, -18, 39, -29, -21, 1),
                (0, 0, 0, 0, 0, 0, 0, 1, -4, 43, -14, -17, -53, -46, -4),
                (0, 0, 0, 0, 0, 0, 0, -43, 55, -65, 33, -1, 4, -3, -35),
                (0, 0, 0, 0, 0, 0, 0, -34, -3, -13, 10, 44, 1, -6, 5),
                (0, 0, 0, 0, 0, 0, 0, 106, 15, 11, -6, 3, -6, -39, -20),
                (0, 0, 0, 0, 0, 0, 0, -19, 17, 8, -11, 9, -2, -5, 9),
                (0, 0, 0, 0, 0, 0, 0, -8, 47, -2, 2, -41, -14, 117, 15),
                (0, 0, 0, 0, 0, 0, 0, -5, 3, 4, -22, -10, 47, -38, 0),
                (0, 0, 0, 0, 0, 0, 0, -8, 8, 33, 7, 14, 1, -25, -1),
                (0, 0, 0, 0, 0, 0, 0, -2, 4, 12, -2, 5, -41, 20, -27),
                (0, 0, 0, 0, 0, 0, 0, 43, -23, -2, 4, -15, 11, -11, 2),
                (0, 0, 0, 0, 0, 0, 0, 0, -18, -21, 4, 25, -5, -169, 0),
                (0, 0, 0, 0, 0, 0, 0, 15, -1, 1, -4, -32, -12, 11, -18),
                (0, 0, 0, 0, 0, 0, 0, -22, 11, 25, 3, -1, 4, -4, 13),
                (0, 0, 0, 0, 0, 0, 0, 15, 98, 36, -9, 2, -10, -27, 2),
                (0, 0, 0, 0, 0, 0, 0, 3, -10, 17, -22, 15, -1, 18, -16),
                (0, 0, 0, 0, 0, 0, 0, 0, -61, 21, -44, 0, 10, -1, -16),
                (0, 0, 0, 0, 0, 0, 0, -17, 26, -28, 37, -13, 9, 5, -5),
                (0, 0, 0, 0, 0, 0, 0, 33, -8, -29, 2, 27, 1, -28, -3),
                (0, 0, 0, 0, 0, 0, 0, 2, -19, -4, 19, 25, -9, 4, -1),
                (0, 0, 0, 0, 0, 0, 0, 30, 3, 3, -23, -10, 1, -5, 6),
                (0, 0, 0, 0, 0, 0, 0, -49, -4, 1, -3, 58, -15, 16, 1),
                (0, 0, 0, 0, 0, 0, 0, -19, 32, -6, -28, -1, 5, 3, -11),
                (0, 0, 0, 0, 0, 0, 0, 0, 8, -7, 0, 20, -39, -9, 34),
                (0, 0, 0, 0, 0, 0, 0, -15, 8, -3, 2, 14, 1, -2, -30),
                (0, 0, 0, 0, 0, 0, 0, -12, 18, -20, 15, 3, -3, -3, 2),
                (0, 0, 0, 0, 0, 0, 0, 33, -20, -11, 26, -22, 6, -1, 3),
                (0, 0, 0, 0, 0, 0, 0, 28, 1, -17, 0, -39, 5, 5, -29),
                (0, 0, 0, 0, 0, 0, 0, -3, 10, 2, -4, -1, -15, 4, -9),
                (0, 0, 0, 0, 0, 0, 0, 33, -13, 0, -17, 4, 18, -1, -42),
                (0, 0, 0, 0, 0, 0, 0, 13, -19, -112, 3, 1, -2, -1, 13),
                (0, 0, 0, 0, 0, 0, 0, 46, 5, 33, 0, -45, -2, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, 6, -8, -14, -2, 14, 1, -1, 2),
                (0, 0, 0, 0, 0, 0, 0, 31, -17, 2, -5, 7, -7, -16, 1),
                (0, 0, 0, 0, 0, 0, 0, 0, -8, -52, 28, 6, 41, -28, 3),
                (0, 0, 0, 0, -148, 0, 0, -54, 15, -25, 18, -29, 0, -148, -148),
                (0, 0, 0, 0, 0, 0, 0, 0, -46, 3, 44, -23, 0, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, 7, 0, 10, -20, -16, 5, -46, -9),
                (0, 0, 0, 0, 0, 0, 0, 12, 0, 0, -23, -19, -1, 16, 1),
                (0, 0, 0, 0, 0, 0, 0, 39, -19, -2, 2, -15, 15, 4, -2),
                (0, 0, 0, 0, 0, 0, 0, -4, 0, -2, 12, 10, -5, -33, 0),
                (0, 0, 0, 0, 0, 0, 0, -4, 1, 2, -18, -34, 27, 11, -5),
                (0, 0, 0, 0, 0, 0, 0, -4, 2, -36, 4, 8, -8, -10, 10),
                (0, 0, 0, 0, 0, 0, 0, -8, 48, -29, -4, 2, -4, 9, 0),
                (0, 0, 0, 0, 0, 0, 0, -23, 56, 42, -7, -2, 4, 4, -2),
                (0, 0, 0, 0, 0, 0, 0, 30, 4, -1, -23, -16, 1, 18, 3),
                (0, 0, 0, 0, 0, 0, 0, 0, -67, 16, 74, 8, -27, -20, 30),
                (0, 0, 0, 0, 0, 0, 0, -6, 0, -3, -36, -6, 73, -34, -1),
                (0, 0, 0, 0, 0, 0, 0, -51, 7, -1, 50, 0, 5, -3, 0),
                (0, 0, 0, 0, 0, 0, 0, -21, 3, 12, -3, 0, 33, 0, -4),
                (0, 0, 0, 0, 0, 0, 0, 1, -15, 11, 144, -1, 15, -6, -1),
                (0, 0, 0, 0, 0, 0, 0, 0, -14, 52, -20, -32, -11, -8, 4),
                (0, 0, 0, 0, 0, 0, 0, 0, 5, -6, 2, -9, 15, 12, -5),
                (0, 0, 0, 0, 0, 0, 0, 5, 45, -2, -20, 50, 8, 0, 2),
                (0, 0, 0, 0, 0, 0, 0, -18, 24, 12, -54, 31, -3, -36, 0),
                (0, 0, 0, 0, 0, 0, 0, -9, 20, 2, -3, -1, -28, 4, -4),
                (0, 0, 0, 0, 0, 0, 0, -8, 21, 9, -12, 8, 73, 0, -1),
                (0, 0, 0, 0, 0, 0, 0, 0, 9, -14, 35, 13, -5, 9, -4),
                (0, 0, 0, 0, 0, 0, 0, 0, -2, 14, -43, 19, 54, 7, -2),
                (0, 0, 0, 0, 0, 0, 0, 18, -46, 61, 0, 22, -97, 0, 1),
                (0, 0, 0, 0, 0, 0, 0, -11, 1, 7, 0, 3, 29, 1, -18),
                (0, 0, 0, 0, 0, 0, 0, 51, 2, -1, 47, -21, 1, 13, 0),
                (0, 0, 0, 0, 0, 0, 0, 0, 8, -9, 0, -10, 3, -3, -18),
                (0, 0, 0, 0, 0, 0, 0, -2, 5, 0, -5, 5, 0, -27, 8),
                (0, 0, 0, 0, 0, 0, 0, -3, 6, 3, -8, 9, -13, 3, -3),
                (0, 0, 0, 0, 0, 0, 0, 0, 38, 0, -73, 4, 33, -14, 29),
                (0, 0, 0, 0, 0, 0, 0, 0, -26, 0, 84, -2, 3, -3, -24),
                (0, 0, 0, 0, 0, 0, 0, 0, 107, 0, -37, 113, -11, -30, 14),
                (0, 0, 0, 0, 0, 0, 0, -21, 4, 44, 7, 22, -45, 0, -14),
                (0, 0, 0, 0, 0, 0, 0, 0, 1, 28, -38, -114, 0, 27, -2),
                (0, 0, 0, 0, 0, 0, 0, -22, 27, -24, 12, 0, -126, 30, 0),
                (0, 0, 0, 0, 0, 0, 0, 7, -6, 0, -26, 1, -4, -1, 2),
                (0, 0, 0, 0, 0, 0, 0, -2, 4, -9, 9, 13, -3, -1, 5),
                (0, 0, 0, 0, 0, 0, 0, -4, 5, 2, -42, 31, 0, 3, -5)
                );
    constant parent : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 6, 6, 5, 5),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 5, 5, 6, 6, 4, 4),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 5, 5, 6, 6, 4, 4),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6)
                );
    constant depth : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3)
                );
    constant iLeaf : intArray2D(nTrees-1 downto 0)(nLeaves-1 downto 0) := ((7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14)
                );
    constant value : tyArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := to_tyArray2D(value_int);
      constant threshold : txArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := to_txArray2D(threshold_int);
end Arrays0;