library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_misc.all;
  use ieee.numeric_std.all;

  use work.Constants.all;
  use work.Types.all;
  package Arrays0 is

    constant initPredict : ty := to_ty(0);
    constant feature : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((4, 1, 0, 3, 1, 0, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 1, 0, 0, 1, 3, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 1, 0, 0, 19, 0, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 4, 4, 3, 1, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 3, 0, 17, 1, 3, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 4, 0, 4, 1, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 1, 3, 4, 0, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 3, 3, 17, 20, 0, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 4, 1, 16, 2, 17, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 4, 2, 3, 17, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 0, 4, 1, 4, 1, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 4, 17, 0, 16, 7, 12, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 16, 18, 12, 1, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 18, 4, 4, 18, 16, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 20, 5, 16, 13, 6, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 7, 4, 17, 6, 20, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 4, 18, 18, 0, 0, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 18, 16, 4, 2, 20, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 7, 16, 17, 6, 1, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 17, 20, 7, 14, 10, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 1, 16, 18, 16, 1, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 4, 18, 16, 0, 5, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 2, 17, 7, 16, 7, 12, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 17, 20, 7, 13, 17, 8, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 17, 20, 7, 18, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 5, 17, 8, 16, 7, 12, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 20, 2, 17, 16, 1, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 18, 16, 18, 2, 2, 15, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 2, 16, 6, 18, 1, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 18, 18, 20, 1, 5, 20, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 17, 8, 6, 19, 17, 5, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 2, 17, -2, 19, 7, 14, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 17, 1, 3, 17, 16, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 3, 17, 17, 16, 2, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 1, 4, 18, 16, 1, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 15, 4, 17, 4, 3, 13, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 20, 16, 17, 16, 0, 5, -2, -2, -2, -2, -2, -2, -2, -2),
                (6, 16, 19, 4, 2, 11, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 17, 1, 17, 0, 5, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 18, 17, 18, 4, 16, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 16, 16, 17, 19, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 4, 4, 16, 16, 0, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 4, 2, 19, 16, 16, 5, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 4, 19, 5, 16, 10, 12, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 16, 16, 4, 5, 17, 10, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 17, 1, 19, 14, 16, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (15, 17, 13, 13, 14, 17, 14, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 4, 18, 16, 16, 4, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (6, 17, 16, 4, 19, 4, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 20, 17, 10, 2, 7, 12, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 2, 19, 18, 17, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 16, 4, 4, 4, 0, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 2, 0, -2, 17, 16, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (6, 16, 17, 4, 2, 0, 9, -2, -2, -2, -2, -2, -2, -2, -2),
                (19, 5, 12, 7, 7, 15, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (15, 20, 17, 17, 13, 12, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 8, 17, 0, 5, 5, 10, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 19, 15, 4, 3, 17, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 16, 17, 0, 2, 16, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 18, 16, 4, 18, 19, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 4, 19, 10, 10, 11, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 6, 3, 16, 3, 2, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 16, 16, 4, 4, 4, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 18, 17, 0, 3, 16, 6, -2, -2, -2, -2, -2, -2, -2, -2),
                (7, 13, 13, 10, 12, 17, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (10, 1, 4, 17, 3, 7, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 0, 2, 1, 16, 1, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 5, 18, 17, 16, 20, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (7, 13, 13, 10, 12, 17, 11, -2, -2, -2, -2, -2, -2, -2, -2),
                (10, 4, 4, 16, 17, 7, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (7, 13, 13, 10, 3, 10, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 1, 4, 8, 10, 16, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 20, 0, 12, 5, 1, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 1, 3, 16, 16, 16, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 2, 17, 20, 10, 16, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 0, 16, -2, 16, 0, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 20, 15, 17, 17, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 7, 17, 17, 13, 16, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 1, 18, 5, 16, 20, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 17, 4, 17, 16, 17, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 1, 16, 16, 3, 2, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 16, 4, 8, 1, 0, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 0, 18, -2, -2, 4, 14, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 2, 17, 4, 10, 16, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 0, 16, 1, -2, 2, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 16, 1, 9, -2, 16, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 5, 2, 9, 2, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (9, 10, 16, 17, 4, 8, 5, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 20, 3, 20, 17, 12, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 17, 4, 2, 2, 1, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (11, 0, 7, 16, 17, 19, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 2, 1, 4, 3, 14, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 16, 16, 20, 2, 0, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 16, 3, 2, 2, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 17, 9, 5, 9, 16, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 16, 16, 4, 2, 0, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 17, 3, 18, 3, 0, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (19, 17, 4, 20, 12, 2, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (15, 17, 17, 20, 14, 12, 14, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 17, 2, 17, 3, 2, 3, -2, -2, -2, -2, -2, -2, -2, -2)
                );
    constant threshold_int : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((576, 205, 3542, 514, 327, 1723, 978, 0, 0, 0, 0, 0, 0, 0, 0),
                (576, 177, 4115, 2500, 292, 1302, 808, 0, 0, 0, 0, 0, 0, 0, 0),
                (576, 227, 2782, 1037, 320, 1428, 263, 0, 0, 0, 0, 0, 0, 0, 0),
                (280, 2480, 704, 576, 878, 448, 7466, 0, 0, 0, 0, 0, 0, 0, 0),
                (576, 412, 7372, 400, 107, 1201, 1166, 0, 0, 0, 0, 0, 0, 0, 0),
                (312, 1903, 704, 917, 704, 533, 1461, 0, 0, 0, 0, 0, 0, 0, 0),
                (242, 11782, 391, 1058, 576, 1071, 580, 0, 0, 0, 0, 0, 0, 0, 0),
                (704, 629, 1424, 460, 192, 27265, 16914, 0, 0, 0, 0, 0, 0, 0, 0),
                (1326, 576, 372, 299921, 439, 395, 145, 0, 0, 0, 0, 0, 0, 0, 0),
                (152, 1591, 704, 275, 1292, 126, 13621, 0, 0, 0, 0, 0, 0, 0, 0),
                (709, 23908, 704, 492, 576, 122, 1519, 0, 0, 0, 0, 0, 0, 0, 0),
                (1148, 576, 415, 498, 192686, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (526, 8525, 309262, 1241, 64, 687, 263, 0, 0, 0, 0, 0, 0, 0, 0),
                (738, -1166, 576, 704, 1084, 252138, 19261, 0, 0, 0, 0, 0, 0, 0, 0),
                (137, 47508, 192, 64, 29776, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (734, 64, 704, 285, 64, 192, 176196, 0, 0, 0, 0, 0, 0, 0, 0),
                (-979, 576, 1234, -1354, 1646, 40262, 576, 0, 0, 0, 0, 0, 0, 0, 0),
                (1379, -1339, 208063, 576, 236, 576, 370231, 0, 0, 0, 0, 0, 0, 0, 0),
                (645, 64, 308622, 285, 64, 796, 485, 0, 0, 0, 0, 0, 0, 0, 0),
                (578, 549, 576, 64, 64, 64, 12252, 0, 0, 0, 0, 0, 0, 0, 0),
                (47835, 761, 27652, 1414, 316378, 31, 149, 0, 0, 0, 0, 0, 0, 0, 0),
                (-896, 576, 739, 375762, 1609, 64, 576, 0, 0, 0, 0, 0, 0, 0, 0),
                (705, 109, 270, 64, 51223, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (950, 382, 576, 64, 64, 101, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (352, 116, 576, 64, 986, 113777, 223542, 0, 0, 0, 0, 0, 0, 0, 0),
                (66, 64, 284, 64, 236120, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (195, 576, 57284, 81, 297291, 888, 18176, 0, 0, 0, 0, 0, 0, 0, 0),
                (1644, -1354, 208063, -1669, 35665, 6438, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (645, 70, 292840, 64, 1534, 916, 373772, 0, 0, 0, 0, 0, 0, 0, 0),
                (-731, -1541, 656, 576, 107, 64, 576, 0, 0, 0, 0, 0, 0, 0, 0),
                (469, 105, 64, 64, 192, 280, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (3035, 1686, 293, 0, 448, 64, 64, 0, 0, 0, 0, 0, 0, -256, -256),
                (321, 30, 97, 183, 188, 301237, 262, 0, 0, 0, 0, 0, 0, 0, 0),
                (72002, 1644, 249, 555, 229409, 84108, 39589, 0, 0, 0, 0, 0, 0, 0, 0),
                (382944, 916, 576, -656, 376335, 236, -4, 0, 0, 0, 0, 0, 0, 0, 0),
                (1549, 64, 704, 376, 576, 4228, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (438, 576, 4350, 102, 231298, 3053, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (64, 140417, 192, 576, 2331, 64, 246, 0, 0, 0, 0, 0, 0, 0, 0),
                (70, 196, 64, 122, 203, 64, 121, 0, 0, 0, 0, 0, 0, 0, 0),
                (4123, 1639, 638, -1661, 704, 363318, 576, 0, 0, 0, 0, 0, 0, 0, 0),
                (955, 65938, 270550, 3035, 142, 320, 376335, 0, 0, 0, 0, 0, 0, 0, 0),
                (381461, 704, 576, 134111, 223643, 14795, 266, 0, 0, 0, 0, 0, 0, 0, 0),
                (-1339, 576, 438, 320, 106460, 51527, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (74, 704, 192, 64, 140991, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (13949, 44310, 24347, 576, 64, 396, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (74, 246, 39, 192, 64, 228971, 814, 0, 0, 0, 0, 0, 0, 0, 0),
                (64, 384, 64, 64, 64, 405, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (-566, 576, 619, 179029, 254363, 576, 704, 0, 0, 0, 0, 0, 0, 0, 0),
                (64, 137, 305620, 576, 448, 704, 576, 0, 0, 0, 0, 0, 0, 0, 0),
                (140, 576, 254, 64, 38, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (2102, 84960, 576, 1414, 200, 235412, 378830, 0, 0, 0, 0, 0, 0, 0, 0),
                (378459, 327776, 576, 576, 576, 13361, 1308, 0, 0, 0, 0, 0, 0, 0, 0),
                (3035, 2211, 1609, 0, 170, 47143, 248, 0, 0, 0, 0, 0, 0, -256, -256),
                (64, 109899, 186, 576, 3971, 5068, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (192, 64, 64, 64, 64, 64, 303, 0, 0, 0, 0, 0, 0, 0, 0),
                (64, 192, 355, 265, 64, 64, 576, 0, 0, 0, 0, 0, 0, 0, 0),
                (105, 64, 177, 2479, 64, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (-1661, 320, 64, 576, 302, 376, 369, 0, 0, 0, 0, 0, 0, 0, 0),
                (985, 5429, 251, 3090, 47, 316445, 500, 0, 0, 0, 0, 0, 0, 0, 0),
                (2376, -566, 369490, 704, 619, 576, 371985, 0, 0, 0, 0, 0, 0, 0, 0),
                (58, 576, 192, 64, 64, 64, 241, 0, 0, 0, 0, 0, 0, 0, 0),
                (118724, 64, 649, 183615, 4137, 121978, 819, 0, 0, 0, 0, 0, 0, 0, 0),
                (263, 260602, 187729, 576, 576, 576, 253, 0, 0, 0, 0, 0, 0, 0, 0),
                (1145, 1714, 148, 79187, 885, 338263, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (64, 64, 64, 64, 64, 249, 576, 0, 0, 0, 0, 0, 0, 0, 0),
                (64, 281, 576, 127, 399, 64, 124568, 0, 0, 0, 0, 0, 0, 0, 0),
                (383417, 277, 18052, 582, 6677, 186, 0, 0, 0, 0, 0, 0, 0, -256, -256),
                (41, 64, -1721, 180, 160684, 192, 54, 0, 0, 0, 0, 0, 0, 0, 0),
                (64, 64, 64, 64, 64, 265, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (64, 576, 576, 142373, 127, 64, 4970, 0, 0, 0, 0, 0, 0, 0, 0),
                (64, 64, 64, 64, 660, 64, 576, 0, 0, 0, 0, 0, 0, 0, 0),
                (326629, 670, 576, 64, 64, 369523, 494, 0, 0, 0, 0, 0, 0, 0, 0),
                (732, 64, 11021, 64, 64, 127, 0, 0, 0, 0, 0, 0, 0, -256, -256),
                (107413, 278, 648, 260939, 260467, 18007, 810, 0, 0, 0, 0, 0, 0, 0, 0),
                (1145, 69, 266, 576, 64, 339207, 400, 0, 0, 0, 0, 0, 0, 0, 0),
                (68, 28, 3035, 0, 359643, 4320, 18480, 0, 0, 0, 0, 0, 0, -256, -256),
                (735, 64, 64, 573, 308, 0, 0, 0, 0, 0, 0, -256, -256, -256, -256),
                (80483, 64, 608, 297, 64, 79111, 495, 0, 0, 0, 0, 0, 0, 0, 0),
                (41, 41, -1744, 64, 74019, 192, 23, 0, 0, 0, 0, 0, 0, 0, 0),
                (1706, 419, 704, 308, 69905, 466, 0, 0, 0, 0, 0, 0, 0, -256, -256),
                (601, 280, 344738, 328012, 884, 5369, -769, 0, 0, 0, 0, 0, 0, 0, 0),
                (371310, 351145, 576, 64, 301, 26090, 1045, 0, 0, 0, 0, 0, 0, 0, 0),
                (2394, 4400, -566, 0, 0, 576, 64, 0, 0, 0, 0, -256, -256, -256, -256),
                (1145, 285, 168, 576, 64, 340050, 123, 0, 0, 0, 0, 0, 0, 0, 0),
                (11, 905, 384057, 407, 0, 2554, 2987, 0, 0, 0, 0, 0, 0, -256, -256),
                (68, 360385, 104, 64, 0, 171678, 806, 0, 0, 0, 0, 0, 0, -256, -256),
                (187, 64, 2554, 64, 1892, 63667, 69669, 0, 0, 0, 0, 0, 0, 0, 0),
                (64, 64, 151445, 206, 576, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (262, 320, 657, 192, 219, 64, 557, 0, 0, 0, 0, 0, 0, 0, 0),
                (370096, 187, 576, 5006, 3695, 242, -431, 0, 0, 0, 0, 0, 0, 0, 0),
                (64, 1488, 64, 32373, 321, 320, 576, 0, 0, 0, 0, 0, 0, 0, 0),
                (6980, 3413, 19, 576, 849, 64, 20, 0, 0, 0, 0, 0, 0, 0, 0),
                (704, 87373, 135663, 576, 2044, 7229, 557, 0, 0, 0, 0, 0, 0, 0, 0),
                (735, 6340, 1179, 3511, 10, 0, 0, 0, 0, 0, 0, -256, -256, -256, -256),
                (187, 138, 64, 64, 64, 207794, 4463, 0, 0, 0, 0, 0, 0, 0, 0),
                (704, 87373, 150669, 576, 1425, 3333, 439, 0, 0, 0, 0, 0, 0, 0, 0),
                (277, 49, 5, -514, 5, 1840, 704, 0, 0, 0, 0, 0, 0, 0, 0),
                (448, 314, 704, 320, 64, 273, 1091, 0, 0, 0, 0, 0, 0, 0, 0),
                (64, 376, 345, 192, 64, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (671, 670, 20381, 424, 517, 17604, 656, 0, 0, 0, 0, 0, 0, 0, 0)
                );
    constant children_left : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 13, 7, 9, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 13, 7, 9, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 13, 7, 9, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 11, 13, 7, 9, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 13, 9, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 13, 9, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1)
                );
    constant children_right : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 14, 8, 10, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 14, 8, 10, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 14, 8, 10, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 12, 14, 8, 10, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 14, 10, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 14, 10, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1)
                );
    constant value_int : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((0, 0, 0, 0, 0, 0, 0, 9, -42, -45, -62, 61, 43, 11, -47),
                (0, 0, 0, 0, 0, 0, 0, 28, -21, -31, -49, 46, -25, 9, -33),
                (0, 0, 0, 0, 0, 0, 0, 34, -16, -42, -20, 42, 29, 8, -33),
                (0, 0, 0, 0, 0, 0, 0, 15, 36, 5, -29, -27, -40, 28, -16),
                (0, 0, 0, 0, 0, 0, 0, -15, 36, -13, -35, 29, -18, -1, -31),
                (0, 0, 0, 0, 0, 0, 0, 32, 20, -10, 15, -23, -36, 29, -7),
                (0, 0, 0, 0, 0, 0, 0, 20, -18, -22, -5, 22, -14, -22, -34),
                (0, 0, 0, 0, 0, 0, 0, -4, 31, -8, -28, 23, -6, -15, -32),
                (0, 0, 0, 0, 0, 0, 0, -9, 19, 29, 19, -6, 14, -32, -19),
                (0, 0, 0, 0, 0, 0, 0, 27, 17, 7, -17, -26, -7, 15, -7),
                (0, 0, 0, 0, 0, 0, 0, 11, -19, -24, -5, -9, -24, 7, -19),
                (0, 0, 0, 0, 0, 0, 0, 20, -6, 29, 18, -20, -2, -28, 14),
                (0, 0, 0, 0, 0, 0, 0, 8, -29, -14, 0, -19, -31, 16, -10),
                (0, 0, 0, 0, 0, 0, 0, -31, 13, 7, -21, -25, -10, 1, -16),
                (0, 0, 0, 0, 0, 0, 0, 19, 5, -32, -13, -22, 14, -27, -6),
                (0, 0, 0, 0, 0, 0, 0, -29, 17, -15, 24, 9, -9, 16, -3),
                (0, 0, 0, 0, 0, 0, 0, -33, -19, 12, -8, 4, -14, -30, -2),
                (0, 0, 0, 0, 0, 0, 0, -30, -13, 16, 1, -24, -11, -11, 10),
                (0, 0, 0, 0, 0, 0, 0, -33, 5, -19, 7, -19, -29, 10, -12),
                (0, 0, 0, 0, 0, 0, 0, -5, 6, 34, 10, -8, -24, 9, -9),
                (0, 0, 0, 0, 0, 0, 0, 2, -23, -27, -2, 3, -32, -7, -17),
                (0, 0, 0, 0, 0, 0, 0, -19, 14, 10, -6, 11, 1, -15, 1),
                (0, 0, 0, 0, 0, 0, 0, 11, 24, 30, 4, -29, 0, -19, 6),
                (0, 0, 0, 0, 0, 0, 0, -11, 3, -23, 11, -21, -8, -26, 1),
                (0, 0, 0, 0, 0, 0, 0, -24, -1, 7, -8, -13, -3, 9, -5),
                (0, 0, 0, 0, 0, 0, 0, 8, 36, 8, 0, -22, -1, -16, 5),
                (0, 0, 0, 0, 0, 0, 0, -12, 11, 24, 13, 0, -24, -35, -12),
                (0, 0, 0, 0, 0, 0, 0, -29, -13, 2, -7, -21, -14, 1, -15),
                (0, 0, 0, 0, 0, 0, 0, -1, 19, 0, -19, -14, -27, -1, 32),
                (0, 0, 0, 0, 0, 0, 0, -21, -1, 0, -7, 8, 1, -7, 5),
                (0, 0, 0, 0, 0, 0, 0, -28, -1, 9, 2, -12, -2, 19, -2),
                (0, 0, 0, -11, 0, 0, 0, -43, -71, -17, 1, 12, -1, -11, -11),
                (0, 0, 0, 0, 0, 0, 0, -15, 19, 20, 9, 5, -2, -4, 1),
                (0, 0, 0, 0, 0, 0, 0, 0, 8, -13, -2, -11, -22, -31, -5),
                (0, 0, 0, 0, 0, 0, 0, -4, 1, -21, 35, 29, 59, 8, -19),
                (0, 0, 0, 0, 0, 0, 0, -1, 12, -19, 0, -21, 17, 34, 3),
                (0, 0, 0, 0, 0, 0, 0, -10, 4, 21, 7, 4, -41, 3, -2),
                (0, 0, 0, 0, 0, 0, 0, -25, -5, -8, 6, 2, 28, -12, 0),
                (0, 0, 0, 0, 0, 0, 0, 10, 28, 14, -6, 12, 2, 3, -2),
                (0, 0, 0, 0, 0, 0, 0, -19, 0, -21, 17, -15, 7, 22, -11),
                (0, 0, 0, 0, 0, 0, 0, -36, 0, -17, -6, -29, -6, -9, 22),
                (0, 0, 0, 0, 0, 0, 0, -8, 1, 9, -8, 29, -12, -1, -22),
                (0, 0, 0, 0, 0, 0, 0, -16, -2, 13, -6, 24, 3, 3, -1),
                (0, 0, 0, 0, 0, 0, 0, 11, -13, 16, -5, 8, -3, -14, 0),
                (0, 0, 0, 0, 0, 0, 0, -20, 23, 4, -1, -21, -46, 1, -9),
                (0, 0, 0, 0, 0, 0, 0, 2, -16, 21, 1, 8, 1, -1, -12),
                (0, 0, 0, 0, 0, 0, 0, 1, -7, 29, -1, -4, -29, -15, 2),
                (0, 0, 0, 0, 0, 0, 0, -14, -1, 4, -6, 4, 0, -5, 4),
                (0, 0, 0, 0, 0, 0, 0, -23, 10, 7, -4, 0, 5, 8, -9),
                (0, 0, 0, 0, 0, 0, 0, 4, -16, 24, 13, -13, 0, -7, 2),
                (0, 0, 0, 0, 0, 0, 0, 1, -9, -17, -6, -9, 3, -20, 5),
                (0, 0, 0, 0, 0, 0, 0, -2, 2, 5, -8, 19, -9, -8, 22),
                (0, 0, 0, -3, 0, 0, 0, -29, -41, 24, 0, -2, 1, -3, -3),
                (0, 0, 0, 0, 0, 0, 0, -20, -6, -5, 5, 6, -3, 0, -11),
                (0, 0, 0, 0, 0, 0, 0, 80, 5, -15, 2, -17, 9, -4, 2),
                (0, 0, 0, 0, 0, 0, 0, 75, 7, 1, -3, 36, 8, -17, -2),
                (0, 0, 0, 0, 0, 0, 0, -4, -23, 9, -3, 20, 3, 0, -11),
                (0, 0, 0, 0, 0, 0, 0, -23, -3, 19, -14, 0, 6, 10, -4),
                (0, 0, 0, 0, 0, 0, 0, 9, -33, 8, 0, -27, -3, 5, -18),
                (0, 0, 0, 0, 0, 0, 0, -3, 2, 1, -2, -4, -16, 42, 6),
                (0, 0, 0, 0, 0, 0, 0, -2, -19, -17, 3, 1, 16, -6, 0),
                (0, 0, 0, 0, 0, 0, 0, -8, 1, 1, -14, -26, -1, -48, -13),
                (0, 0, 0, 0, 0, 0, 0, -4, 3, 3, -6, -8, 1, 12, 2),
                (0, 0, 0, 0, 0, 0, 0, 0, -6, -18, 7, -30, -11, -27, -3),
                (0, 0, 0, 0, 0, 0, 0, -14, 6, -8, 3, 1, 16, -28, -2),
                (0, 0, 0, 0, 0, 0, 0, -5, 0, 7, -1, 7, -27, 8, -3),
                (0, 0, 0, 0, 0, 0, -24, 8, -17, -13, 0, 7, 24, -24, -24),
                (0, 0, 0, 0, 0, 0, 0, 23, 3, 6, 0, 6, -19, 3, 0),
                (0, 0, 0, 0, 0, 0, 0, -11, 3, -6, 2, 1, 14, -21, 0),
                (0, 0, 0, 0, 0, 0, 0, -7, 5, -13, 0, 3, -23, 5, -6),
                (0, 0, 0, 0, 0, 0, 0, -9, 1, 2, -3, 4, -2, -21, 0),
                (0, 0, 0, 0, 0, 0, 0, 0, 2, -5, -18, 0, 11, 3, -7),
                (0, 0, 0, 0, 0, 0, 3, 23, -6, 2, 0, 24, 52, 3, 3),
                (0, 0, 0, 0, 0, 0, 0, 1, -2, -1, 5, -29, -1, -37, -11),
                (0, 0, 0, 0, 0, 0, 0, 2, 16, 0, -1, -25, -5, 9, -23),
                (0, 0, 0, -10, 0, 0, 0, 34, 10, -1, -33, 5, 0, -10, -10),
                (0, 0, 0, 0, 0, 7, 40, -12, 0, 0, 1, 7, 7, 40, 40),
                (0, 0, 0, 0, 0, 0, 0, -6, 0, 1, -2, -9, 0, -46, -16),
                (0, 0, 0, 0, 0, 0, 0, 7, 1, -8, 22, 5, -18, -3, 0),
                (0, 0, 0, 0, 0, 0, 22, 0, 3, -11, -1, -17, 10, 22, 22),
                (0, 0, 0, 0, 0, 0, 0, 0, -2, 3, -3, -10, 0, -18, 11),
                (0, 0, 0, 0, 0, 0, 0, -1, 1, -4, 6, 9, -25, -4, 9),
                (0, 0, 0, -17, -31, 0, 0, -3, 0, 1, -1, -17, -17, -31, -31),
                (0, 0, 0, 0, 0, 0, 0, -4, 7, 0, -2, -28, -5, 20, -13),
                (0, 0, 0, 0, -8, 0, 0, 17, -5, -1, 0, 18, -7, -8, -8),
                (0, 0, 0, 0, -11, 0, 0, 37, 10, 3, 0, 0, -3, -11, -11),
                (0, 0, 0, 0, 0, 0, 0, -20, 12, 3, -3, 18, -5, -10, 2),
                (0, 0, 0, 0, 0, 0, 0, 10, 0, -20, 8, -12, 5, 11, -6),
                (0, 0, 0, 0, 0, 0, 0, 41, -13, 0, 4, -4, 2, -4, 2),
                (0, 0, 0, 0, 0, 0, 0, 2, -2, -3, 1, 4, 14, 6, -4),
                (0, 0, 0, 0, 0, 0, 0, 24, 0, -2, 1, -10, 0, 7, 1),
                (0, 0, 0, 0, 0, 0, 0, -24, 28, -34, -6, 8, -6, -26, 0),
                (0, 0, 0, 0, 0, 0, 0, -9, 2, -3, 2, 17, 0, 6, -3),
                (0, 0, 0, 0, 0, 35, 0, 7, -25, 11, 0, 35, 35, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, 6, -2, 14, 3, -2, 1, -12, -3),
                (0, 0, 0, 0, 0, 0, 0, -8, 0, -3, 2, 16, 1, 6, -2),
                (0, 0, 0, 0, 0, 0, 0, -34, -3, -29, 8, -3, 16, 0, 1),
                (0, 0, 0, 0, 0, 0, 0, -4, 0, -6, 5, 11, -5, 0, 14),
                (0, 0, 0, 0, 0, 0, 0, 8, 0, 14, -3, 30, 4, -12, -1),
                (0, 0, 0, 0, 0, 0, 0, 0, -1, -53, -9, 7, 34, -35, 1)
                );
    constant parent : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 4, 4, 5, 5, 6, 6, 3, 3),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 4, 4, 5, 5, 6, 6, 3, 3),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 4, 4, 5, 5, 6, 6, 3, 3),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 5, 5, 6, 6, 3, 3, 4, 4),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 5, 5, 6, 6, 4, 4),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 5, 5, 6, 6, 4, 4),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6)
                );
    constant depth : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3)
                );
    constant iLeaf : intArray2D(nTrees-1 downto 0)(nLeaves-1 downto 0) := ((7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14)
                );
    constant value : tyArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := to_tyArray2D(value_int);
      constant threshold : txArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := to_txArray2D(threshold_int);
end Arrays0;