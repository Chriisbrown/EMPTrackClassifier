library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_misc.all;
  use ieee.numeric_std.all;

  use work.Constants.all;
  use work.Types.all;
  package Arrays0 is

    constant initPredict : ty := to_ty(0);
    constant feature : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((1, 0, 4, 4, 4, 19, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 4, 4, 3, 1, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 1, 0, 0, 17, 2, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 1, 0, 16, 3, 2, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 4, 4, 4, 16, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 3, 0, 17, 19, 0, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 1, 1, 4, 4, 4, 12, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 1, 1, 4, 4, 4, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 1, 1, 18, 4, 3, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 2, 4, 4, 17, 1, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 16, 0, 10, 18, 0, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 16, 18, 18, 1, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 20, 2, 13, 7, 16, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 18, 4, 4, 18, 1, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 1, 1, 2, 17, 5, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 16, 18, 18, 1, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 17, 2, 5, 16, 16, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 1, 18, 2, 0, 18, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 18, 4, 4, 0, 19, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 7, 3, 17, 6, 12, 14, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 2, 1, 6, 1, 17, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 17, 20, 7, 14, 16, 7, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 18, 16, 5, 16, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 4, 18, 19, 0, 3, 20, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 7, 12, 5, 6, 5, 15, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 16, 17, 17, 17, 7, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 20, 4, 10, 2, 1, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 3, 18, 4, 1, 16, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 7, 16, 12, 13, 10, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 17, 8, 7, 12, 17, 5, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 6, 17, 17, 2, 7, 12, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 1, 0, 5, 19, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 1, 4, 16, 16, 1, 20, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 16, 16, 20, 1, 2, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 6, 18, 17, 17, 16, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 18, 0, 19, 16, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 20, 14, 0, 5, 15, 13, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 4, 17, 5, 16, 17, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 17, 1, 19, 14, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 3, 16, 7, 20, 4, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 16, 2, 17, 2, 0, 5, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 18, 4, 20, 1, 18, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 17, 16, 5, 3, 3, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 4, 19, 6, 2, 10, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 2, 18, 4, 20, 18, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 16, 4, 2, 4, 20, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 1, 10, 19, 4, 6, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (7, 13, 13, 10, 12, 10, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 17, 17, 5, 17, 4, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 1, 16, 1, 16, 2, 19, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 0, 7, 4, 17, 13, 13, -2, -2, -2, -2, -2, -2, -2, -2),
                (6, 16, 17, 20, 2, 5, 10, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 17, 4, 18, 1, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 17, 8, 7, 14, 10, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 16, 0, 1, 6, 5, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 4, 3, 3, 3, 18, 19, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 17, 0, 8, 17, 4, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 6, 14, 20, 0, 12, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 7, 14, 5, 13, 15, 19, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 4, 17, 10, 10, 5, 10, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 4, 18, 2, 2, 4, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 0, 2, -2, -2, 5, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 17, 4, 20, 19, 0, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 19, 19, 16, 2, 14, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 6, 16, 0, 3, 2, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 13, 14, 5, 4, 15, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 9, 2, 10, 16, 4, 8, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 16, 2, 17, 5, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 16, 16, 8, 4, 16, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 18, 17, -2, 3, 20, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 19, 4, 13, 17, 10, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 2, 17, 0, 5, 16, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 2, 14, 12, 16, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (6, 16, 0, 4, 0, 3, 5, -2, -2, -2, -2, -2, -2, -2, -2),
                (19, 11, 17, 8, 1, 0, 12, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 4, 2, 3, 3, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 1, 10, 2, 15, 12, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 16, 3, 0, 20, 1, 7, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 16, 4, 4, 4, 1, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 7, 14, 5, 11, 15, 19, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 17, 9, 6, 2, 19, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 1, 4, 4, 2, 17, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 13, 13, 17, 4, 5, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (8, 10, 5, 16, 2, 7, 7, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 17, 17, 19, -2, 18, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 17, 9, 3, 2, 17, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 3, 17, 3, 0, 17, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 1, 18, 19, 17, -2, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 3, 0, 17, 19, 12, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 20, 6, 16, 11, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 8, 16, -2, 3, 4, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 3, 13, 18, 18, 3, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 12, 1, 3, 11, 19, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 17, 2, 16, 0, 18, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 1, 17, 5, 16, 1, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 20, 18, 19, 1, 5, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 1, 16, 16, -2, 6, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 18, 16, 0, 3, 2, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (5, 2, 2, 16, 17, 4, 9, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 4, 1, 4, 3, 0, -2, -2, -2, -2, -2, -2, -2, -2)
                );
    constant threshold_int : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((304, 2780, 576, 576, 576, 320, 2064, 0, 0, 0, 0, 0, 0, 0, 0),
                (288, 2046, 576, 576, 1166, 516, 2642, 0, 0, 0, 0, 0, 0, 0, 0),
                (576, 190, 3018, 2482, 408, 2046, 3578, 0, 0, 0, 0, 0, 0, 0, 0),
                (576, 226, 2914, 172, 422, 2046, 3336, 0, 0, 0, 0, 0, 0, 0, 0),
                (362, 1996, 704, 576, 704, 272, 2844, 0, 0, 0, 0, 0, 0, 0, 0),
                (576, 540, 2066, 396, 320, 1324, 1216, 0, 0, 0, 0, 0, 0, 0, 0),
                (1650, 572, 204, 576, 576, 704, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (1492, 396, 454, 576, 576, 704, 666, 0, 0, 0, 0, 0, 0, 0, 0),
                (1384, 250, 152, 1294, 576, 1056, 394, 0, 0, 0, 0, 0, 0, 0, 0),
                (882, 2046, 704, 576, 448, 124, 1512, 0, 0, 0, 0, 0, 0, 0, 0),
                (576, 212, 2168, 64, -1136, 922, 872, 0, 0, 0, 0, 0, 0, 0, 0),
                (532, 942, 302, 1421, 1234, 764, 426, 0, 0, 0, 0, 0, 0, 0, 0),
                (704, 192, 2044, 64, 64, 186, 3696, 0, 0, 0, 0, 0, 0, 0, 0),
                (660, -1151, 704, 704, 1091, 104, 1384, 0, 0, 0, 0, 0, 0, 0, 0),
                (732, 228, 122, 194, 120, 64, 278, 0, 0, 0, 0, 0, 0, 0, 0),
                (602, 2396, 336, -1316, -1016, 916, -746, 0, 0, 0, 0, 0, 0, 0, 0),
                (704, 116, 2044, 64, 138, 184, 134, 0, 0, 0, 0, 0, 0, 0, 0),
                (716, 136, 1391, 142, 458, -941, 704, 0, 0, 0, 0, 0, 0, 0, 0),
                (806, -731, 576, 576, 2284, 320, 704, 0, 0, 0, 0, 0, 0, 0, 0),
                (556, 64, 1072, 294, 64, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (560, 70, 764, 64, 202, 390, 356, 0, 0, 0, 0, 0, 0, 0, 0),
                (614, 552, 576, 64, 64, 102, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (104, 1324, 1271, 182, 64, 180, 704, 0, 0, 0, 0, 0, 0, 0, 0),
                (-1338, 576, 731, 320, 1796, 950, 576, 0, 0, 0, 0, 0, 0, 0, 0),
                (384, 64, 64, 64, 64, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (850, 492, 308, 78, 296, 144, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (370, 576, 576, 64, 2046, 300, 1214, 0, 0, 0, 0, 0, 0, 0, 0),
                (-1541, 1948, 1548, 704, 432, 2, 2904, 0, 0, 0, 0, 0, 0, 0, 0),
                (954, 64, 366, 64, 64, 64, 1566, 0, 0, 0, 0, 0, 0, 0, 0),
                (446, 262, 64, 64, 64, 262, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (796, 64, 282, 138, 70, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (2036, 68, 3025, 64, 192, 360, 236, 0, 0, 0, 0, 0, 0, 0, 0),
                (372, 916, 576, 4, 272, 236, 704, 0, 0, 0, 0, 0, 0, 0, 0),
                (-1661, 366, 110, 192, 254, 2046, 1564, 0, 0, 0, 0, 0, 0, 0, 0),
                (284, 64, -566, 626, 190, 364, 626, 0, 0, 0, 0, 0, 0, 0, 0),
                (2036, 1654, 3004, 192, 60, 348, 360, 0, 0, 0, 0, 0, 0, 0, 0),
                (282, 320, 64, 3876, 64, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (74, 704, 184, 64, 170, 136, 246, 0, 0, 0, 0, 0, 0, 0, 0),
                (64, 246, 670, 192, 64, 2, 300, 0, 0, 0, 0, 0, 0, 0, 0),
                (46, 1038, 100, 64, 576, 704, 1564, 0, 0, 0, 0, 0, 0, 0, 0),
                (916, 46, 470, 34, 218, 1264, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (374, -1661, 576, 192, 988, 994, 138, 0, 0, 0, 0, 0, 0, 0, 0),
                (32, 182, 360, 64, 26, 1884, 576, 0, 0, 0, 0, 0, 0, 0, 0),
                (92, 576, 192, 64, 2046, 64, 262, 0, 0, 0, 0, 0, 0, 0, 0),
                (4, 1788, 1721, 576, 704, -566, 614, 0, 0, 0, 0, 0, 0, 0, 0),
                (656, 84, 704, 2044, 576, 576, 2852, 0, 0, 0, 0, 0, 0, 0, 0),
                (990, 300, 64, 320, 576, 64, 216, 0, 0, 0, 0, 0, 0, 0, 0),
                (64, 64, 64, 64, 64, 64, 704, 0, 0, 0, 0, 0, 0, 0, 0),
                (68, 172, 10, 64, 296, 704, 300, 0, 0, 0, 0, 0, 0, 0, 0),
                (640, 300, 284, 246, 138, 2020, 192, 0, 0, 0, 0, 0, 0, 0, 0),
                (2, 2088, 64, 576, 308, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (64, 108, 176, 576, 1166, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (58, 82, 704, -828, 272, 110, 218, 0, 0, 0, 0, 0, 0, 0, 0),
                (462, 246, 64, 64, 64, 64, 186, 0, 0, 0, 0, 0, 0, 0, 0),
                (574, 284, 254, 66, 300, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (-1338, 576, 2036, 1064, 584, 1638, 576, 0, 0, 0, 0, 0, 0, 0, 0),
                (374, 72, 813, 64, 186, 576, 1222, 0, 0, 0, 0, 0, 0, 0, 0),
                (556, 64, 64, 576, 864, 64, 434, 0, 0, 0, 0, 0, 0, 0, 0),
                (312, 64, 64, 64, 64, 64, 320, 0, 0, 0, 0, 0, 0, 0, 0),
                (104, 576, 176, 64, 64, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (-566, 576, 626, 1006, 2006, 576, 576, 0, 0, 0, 0, 0, 0, 0, 0),
                (2, 2088, 46, 0, 0, 64, 1114, 0, 0, 0, 0, -256, -256, -256, -256),
                (370, 686, 576, 64, 448, 774, 2998, 0, 0, 0, 0, 0, 0, 0, 0),
                (32, 448, 320, 224, 382, 64, 240, 0, 0, 0, 0, 0, 0, 0, 0),
                (-1721, 64, 6, 1504, 104, 2039, 1146, 0, 0, 0, 0, 0, 0, 0, 0),
                (324, 64, 64, 64, 704, 64, 342, 0, 0, 0, 0, 0, 0, 0, 0),
                (708, 64, 972, 64, 234, 704, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (1094, 28, 1088, 10, 64, 44, 68, 0, 0, 0, 0, 0, 0, 0, 0),
                (730, 360, 210, 64, 576, 146, 180, 0, 0, 0, 0, 0, 0, 0, 0),
                (66, -854, 644, 0, 6, 64, 390, 0, 0, 0, 0, 0, 0, -256, -256),
                (300, 320, 576, 64, 216, 64, 704, 0, 0, 0, 0, 0, 0, 0, 0),
                (38, 330, 10, 390, 64, 70, 300, 0, 0, 0, 0, 0, 0, 0, 0),
                (916, 44, 64, 64, 6, 284, 278, 0, 0, 0, 0, 0, 0, 0, 0),
                (64, 204, 2448, 576, 2032, 1310, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (192, 64, 240, 64, 306, 3020, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (252, 576, 1114, 406, 1138, 30, 68, 0, 0, 0, 0, 0, 0, 0, 0),
                (532, 300, 64, 200, 64, 64, 704, 0, 0, 0, 0, 0, 0, 0, 0),
                (104, 296, 114, 1532, 576, 298, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (360, 320, 576, 576, 576, 220, 1394, 0, 0, 0, 0, 0, 0, 0, 0),
                (332, 64, 64, 64, 64, 64, 320, 0, 0, 0, 0, 0, 0, 0, 0),
                (186, 134, 64, 64, 140, 192, 224, 0, 0, 0, 0, 0, 0, 0, 0),
                (390, 300, 576, 576, 1150, 458, 3441, 0, 0, 0, 0, 0, 0, 0, 0),
                (308, 64, 64, 262, 576, 64, 580, 0, 0, 0, 0, 0, 0, 0, 0),
                (64, 64, 64, 206, 2046, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (2, 304, 742, 192, 0, 626, 249, 0, 0, 0, 0, 0, 0, -256, -256),
                (186, 136, 64, 356, 188, 206, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (-1661, 1196, 642, 596, 3016, 622, -424, 0, 0, 0, 0, 0, 0, 0, 0),
                (732, 18, -1162, 320, 308, 0, 1184, 0, 0, 0, 0, 0, 0, -256, -256),
                (374, 2036, 2632, 176, 576, 64, 1996, 0, 0, 0, 0, 0, 0, 0, 0),
                (988, 66, 192, 64, 6, 64, 252, 0, 0, 0, 0, 0, 0, 0, 0),
                (2, 64, 34, 0, 526, 576, 1574, 0, 0, 0, 0, 0, 0, -256, -256),
                (1721, 18, 64, -64, -536, 1216, 126, 0, 0, 0, 0, 0, 0, 0, 0),
                (308, 64, 168, 1660, 64, 448, 158, 0, 0, 0, 0, 0, 0, 0, 0),
                (644, 624, 272, 360, 1394, 446, -416, 0, 0, 0, 0, 0, 0, 0, 0),
                (12, 336, 12, 64, 347, 354, 2, 0, 0, 0, 0, 0, 0, 0, 0),
                (-1661, 576, -1654, 320, 142, 64, 734, 0, 0, 0, 0, 0, 0, 0, 0),
                (1214, 1202, 318, 374, 0, 64, 2436, 0, 0, 0, 0, 0, 0, -256, -256),
                (438, 146, 34, 3198, 2038, 2046, 568, 0, 0, 0, 0, 0, 0, 0, 0),
                (64, 1092, 548, 234, 156, 576, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (300, 3192, 576, 254, 704, 1104, 3441, 0, 0, 0, 0, 0, 0, 0, 0)
                );
    constant children_left : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 11, 13, 7, 9, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 13, 7, 9, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 13, 9, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 13, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 13, 7, 9, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 13, 9, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1)
                );
    constant children_right : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 12, 14, 8, 10, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 14, 8, 10, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 14, 10, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 14, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 14, 8, 10, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 14, 10, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1)
                );
    constant value_int : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((0, 0, 0, 0, 0, 0, 0, 24, 61, -37, 9, -57, -27, 60, -9),
                (0, 0, 0, 0, 0, 0, 0, 38, 52, 26, -27, -31, -49, 34, -27),
                (0, 0, 0, 0, 0, 0, 0, 26, -17, -36, 0, 44, 27, -2, -30),
                (0, 0, 0, 0, 0, 0, 0, -16, 21, -12, -36, 40, 22, 5, -21),
                (0, 0, 0, 0, 0, 0, 0, 25, 37, -1, 25, -33, -11, 27, -12),
                (0, 0, 0, 0, 0, 0, 0, -3, 34, -30, -5, 36, 29, 16, -17),
                (0, 0, 0, 0, 0, 0, 0, 21, 33, -27, 20, 4, 21, -25, -3),
                (0, 0, 0, 0, 0, 0, 0, 20, 31, -14, 24, -1, 17, -18, -33),
                (0, 0, 0, 0, 0, 0, 0, 28, -9, -5, 24, 14, -10, -14, 9),
                (0, 0, 0, 0, 0, 0, 0, 8, 27, -3, 25, -6, -24, 11, -20),
                (0, 0, 0, 0, 0, 0, 0, -13, -35, -34, 10, 28, 18, 9, -6),
                (0, 0, 0, 0, 0, 0, 0, 24, -28, 4, -32, -19, -33, 13, -13),
                (0, 0, 0, 0, 0, 0, 0, -19, 20, -23, 2, 31, 18, 9, -17),
                (0, 0, 0, 0, 0, 0, 0, -31, 16, 10, -20, -1, -17, 10, -12),
                (0, 0, 0, 0, 0, 0, 0, 27, 18, -9, 20, 17, 5, -10, 3),
                (0, 0, 0, 0, 0, 0, 0, -27, 9, -21, -2, -18, -32, -22, 14),
                (0, 0, 0, 0, 0, 0, 0, 14, -22, -9, 6, 28, 12, 10, 0),
                (0, 0, 0, 0, 0, 0, 0, 26, 19, 17, 1, -15, 2, -31, 11),
                (0, 0, 0, 0, 0, 0, 0, -15, 2, 9, 0, -23, -4, -5, 10),
                (0, 0, 0, 0, 0, 0, 0, -36, 2, -21, 7, -20, 21, 12, -6),
                (0, 0, 0, 0, 0, 0, 0, 8, 27, 16, 5, -2, 7, -24, 15),
                (0, 0, 0, 0, 0, 0, 0, -6, 6, 29, 11, -18, -6, -31, 6),
                (0, 0, 0, 0, 0, 0, 0, 23, 10, 12, 1, -6, 2, -22, 7),
                (0, 0, 0, 0, 0, 0, 0, -26, -6, 16, -9, 3, -5, -10, 8),
                (0, 0, 0, 0, 0, 0, 0, 20, -19, -16, 5, 4, -36, 20, 0),
                (0, 0, 0, 0, 0, 0, 0, 3, 17, -2, 4, -30, -20, -17, 14),
                (0, 0, 0, 0, 0, 0, 0, 0, -23, 11, 0, 20, 46, -6, 32),
                (0, 0, 0, 0, 0, 0, 0, -25, 15, 12, -22, -51, 1, -24, -4),
                (0, 0, 0, 0, 0, 0, 0, -21, 4, 5, -13, -20, -34, 49, 0),
                (0, 0, 0, 0, 0, 0, 0, -24, 3, -10, 10, -14, -2, 17, -1),
                (0, 0, 0, 0, 0, 0, 0, -25, 5, 22, 7, -19, 0, -14, 4),
                (0, 0, 0, 0, 0, 0, 0, 13, 4, 2, -2, -29, 6, -12, 5),
                (0, 0, 0, 0, 0, 0, 0, -32, 0, -23, -7, 20, 39, 3, -48),
                (0, 0, 0, 0, 0, 0, 0, -8, -25, 0, 46, 14, -8, -3, 3),
                (0, 0, 0, 0, 0, 0, 0, -8, 24, 23, 9, -4, 9, 2, -4),
                (0, 0, 0, 0, 0, 0, 0, 3, -1, 7, -23, -25, -1, -5, 24),
                (0, 0, 0, 0, 0, 0, 0, -16, 80, 12, -1, 14, -10, -17, 2),
                (0, 0, 0, 0, 0, 0, 0, 6, -13, 14, -5, 1, 12, -7, 1),
                (0, 0, 0, 0, 0, 0, 0, 4, -18, 23, 2, -41, 0, -15, 6),
                (0, 0, 0, 0, 0, 0, 0, 7, 21, -24, 17, -9, 8, -3, 2),
                (0, 0, 0, 0, 0, 0, 0, 0, 28, 8, -1, 1, -21, 3, -1),
                (0, 0, 0, 0, 0, 0, 0, -2, -20, 0, -15, 25, -7, 12, -16),
                (0, 0, 0, 0, 0, 0, 0, 28, 10, 24, 1, 0, -6, 14, -5),
                (0, 0, 0, 0, 0, 0, 0, -24, -3, 9, -2, 9, -4, -8, 1),
                (0, 0, 0, 0, 0, 0, 0, -20, 32, -37, 0, -2, 1, -19, 33),
                (0, 0, 0, 0, 0, 0, 0, 13, -7, 4, -1, -6, 3, 8, -11),
                (0, 0, 0, 0, 0, 0, 0, -2, 2, 6, -4, -21, -4, -9, -33),
                (0, 0, 0, 0, 0, 0, 0, -18, 8, -12, 5, 6, -2, -21, 2),
                (0, 0, 0, 0, 0, 0, 0, 21, 4, -3, 3, -13, 2, -1, 2),
                (0, 0, 0, 0, 0, 0, 0, 0, -5, -5, 5, -18, -7, 15, -6),
                (0, 0, 0, 0, 0, 0, 0, -17, 22, -28, -54, -9, 2, 2, -5),
                (0, 0, 0, 0, 0, 0, 0, -17, 7, -10, 3, 10, 1, 0, -16),
                (0, 0, 0, 0, 0, 0, 0, -38, -5, 3, 15, -5, 0, 6, -4),
                (0, 0, 0, 0, 0, 0, 0, -10, 0, 7, 1, -2, -21, 3, -6),
                (0, 0, 0, 0, 0, 0, 0, 29, 8, 0, 2, -16, -5, -9, 6),
                (0, 0, 0, 0, 0, 0, 0, -13, 3, 9, -4, 1, -12, -2, -19),
                (0, 0, 0, 0, 0, 0, 0, -16, -1, 3, 0, 29, 7, 3, 27),
                (0, 0, 0, 0, 0, 0, 0, -7, 12, 4, 0, -32, 14, 12, -1),
                (0, 0, 0, 0, 0, 0, 0, 28, -13, 1, -5, 15, -10, -15, 1),
                (0, 0, 0, 0, 0, 0, 0, -1, -16, -12, 3, 17, 2, 0, -10),
                (0, 0, 0, 0, 0, 0, 0, -10, -2, 6, -2, 3, 0, -4, 1),
                (0, 0, 0, -5, -36, 0, 0, -5, 12, -2, 0, -5, -5, -36, -36),
                (0, 0, 0, 0, 0, 0, 0, -5, 0, 50, 8, 24, 7, -5, 21),
                (0, 0, 0, 0, 0, 0, 0, 10, 1, 18, -8, 0, -12, 3, -4),
                (0, 0, 0, 0, 0, 0, 0, -31, 20, 6, -20, 23, -27, 0, -14),
                (0, 0, 0, 0, 0, 0, 0, 6, -1, -14, 4, 14, -8, 13, -2),
                (0, 0, 0, 0, 0, 0, 0, 2, -14, 2, -6, -12, 4, -2, 3),
                (0, 0, 0, 0, 0, 0, 0, -13, 27, -8, 3, 21, -7, -3, 1),
                (0, 0, 0, 0, 0, 0, 0, -1, 1, 9, -3, 25, -21, 3, 39),
                (0, 0, 0, -2, 0, 0, 0, 8, 35, -5, 0, 6, -9, -2, -2),
                (0, 0, 0, 0, 0, 0, 0, -1, -7, -11, 2, 7, -14, -8, 3),
                (0, 0, 0, 0, 0, 0, 0, -3, 18, 8, 1, -15, -2, 0, 1),
                (0, 0, 0, 0, 0, 0, 0, 12, -5, -9, 0, -20, -2, 27, -7),
                (0, 0, 0, 0, 0, 0, 0, -11, 1, -6, 4, 1, -15, 3, -2),
                (0, 0, 0, 0, 0, 0, 0, -7, 1, 10, 35, -7, 17, -5, 1),
                (0, 0, 0, 0, 0, 0, 0, 2, -12, 11, -12, 22, -3, -2, 1),
                (0, 0, 0, 0, 0, 0, 0, 5, 0, 4, -7, 4, -4, -15, 4),
                (0, 0, 0, 0, 0, 0, 0, 9, 1, 1, -10, -1, 7, -2, 0),
                (0, 0, 0, 0, 0, 0, 0, -1, 1, 2, -5, 3, 13, -4, 14),
                (0, 0, 0, 0, 0, 0, 0, 22, -8, -1, 3, 13, -5, -8, 1),
                (0, 0, 0, 0, 0, 0, 0, -7, 1, 19, 4, 6, -1, -17, -5),
                (0, 0, 0, 0, 0, 0, 0, -1, 1, -5, 5, 2, -9, -9, 11),
                (0, 0, 0, 0, 0, 0, 0, 0, 8, -18, -1, -20, 3, 3, -1),
                (0, 0, 0, 0, 0, 0, 0, -2, 1, -2, -24, 47, 0, -7, 1),
                (0, 0, 0, 0, -39, 0, 0, -15, 12, 0, -1, 7, 39, -39, -39),
                (0, 0, 0, 0, 0, 0, 0, -3, 1, 16, 3, 9, 0, 5, -7),
                (0, 0, 0, 0, 0, 0, 0, -6, -24, 36, -2, 0, -9, -4, 6),
                (0, 0, 0, 0, 0, 37, 0, 9, -5, 0, 1, -9, 32, 37, 37),
                (0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -16, 16, 3, 28, -16),
                (0, 0, 0, 0, 0, 0, 0, -2, 30, -9, 0, 36, -11, 5, -16),
                (0, 0, 0, -32, 0, 0, 0, 1, -23, -15, 9, -2, 0, -32, -32),
                (0, 0, 0, 0, 0, 0, 0, 10, -2, -1, 0, -23, 15, 40, 0),
                (0, 0, 0, 0, 0, 0, 0, 1, -5, -11, -1, 4, 0, 5, -2),
                (0, 0, 0, 0, 0, 0, 0, 0, 2, 12, -8, 22, -1, -5, 4),
                (0, 0, 0, 0, 0, 0, 0, 9, -2, -14, 17, 23, -15, -18, 0),
                (0, 0, 0, 0, 0, 0, 0, -15, 3, 39, 0, -4, 50, 0, 19),
                (0, 0, 0, 0, 34, 0, 0, 0, 8, -30, -9, 19, -14, 34, 34),
                (0, 0, 0, 0, 0, 0, 0, 0, 3, 2, -7, 27, 0, -1, -6),
                (0, 0, 0, 0, 0, 0, 0, -23, -1, 11, 1, -2, 6, 0, -3),
                (0, 0, 0, 0, 0, 0, 0, 0, -4, 7, -6, 5, -7, -4, 9)
                );
    constant parent : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 5, 5, 6, 6, 3, 3, 4, 4),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 4, 4, 5, 5, 6, 6, 3, 3),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 5, 5, 6, 6, 4, 4),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 6, 6, 5, 5),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 4, 4, 5, 5, 6, 6, 3, 3),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 5, 5, 6, 6, 4, 4),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6)
                );
    constant depth : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3)
                );
    constant iLeaf : intArray2D(nTrees-1 downto 0)(nLeaves-1 downto 0) := ((7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14)
                );
    constant value : tyArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := to_tyArray2D(value_int);
      constant threshold : txArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := to_txArray2D(threshold_int);
end Arrays0;