library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_misc.all;
  use ieee.numeric_std.all;

  use work.Constants.all;
  use work.Types.all;
  package Arrays0 is

    constant initPredict : ty := to_ty(0);
    constant feature : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((4, 1, 0, 3, 1, 0, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 1, 0, 0, 17, 3, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 4, 0, 3, 3, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 19, 0, 0, 15, 2, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 1, 3, 0, 3, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 3, 4, 17, 4, 18, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 16, 18, 18, 1, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 17, 5, 16, 4, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 16, 3, 4, 17, 16, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 7, 1, 17, 6, 5, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 0, 4, 3, 2, 5, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (7, 17, 6, 5, 12, 17, 13, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 3, 17, 20, 20, 7, 13, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 17, 1, 7, 14, 0, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 2, 1, 1, 16, 16, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 1, 16, 18, 16, 16, 10, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 10, 4, 1, 4, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 6, 14, 4, 7, 16, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 20, 17, 16, 16, 20, 12, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 1, 17, 3, 16, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 18, 4, 5, 4, 1, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 5, 19, 9, 4, 10, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 2, 1, 4, 3, 5, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 4, 4, 16, 16, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 16, 16, 0, 2, 17, 10, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 17, 3, 17, 13, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 7, 18, 13, 13, 16, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 4, 17, 16, 16, 5, 14, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 4, 4, 8, 2, 18, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 8, 2, 10, 5, 17, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 3, 12, 18, 17, 17, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 7, 14, 10, 11, 15, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 4, 10, 0, 2, 20, 8, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 17, 1, 5, 9, 4, 19, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 18, 16, 19, 4, 19, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 16, 17, 0, 2, 16, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 20, 15, 13, 16, 12, 13, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 2, 17, 4, 16, 5, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 2, 18, 4, 3, 3, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 6, 6, 16, 17, 20, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 17, 0, 16, 16, 17, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 2, 16, -2, 16, 2, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 16, 17, 2, 10, 18, 19, -2, -2, -2, -2, -2, -2, -2, -2),
                (19, 11, 17, 17, 2, 4, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 16, 4, 1, 1, 1, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 3, 19, 9, 4, 16, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (19, 9, 17, 10, 16, 20, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 4, 0, 1, 16, 1, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 13, 1, 5, 3, 4, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 6, 2, 18, 0, 1, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (8, 10, 5, 17, 5, 9, 9, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 18, 6, 17, 17, 0, 20, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 10, 1, 17, 0, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 16, 16, 4, 16, 2, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 17, 17, 4, 2, 2, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 1, 15, 1, 3, 16, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 17, -2, 17, 16, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 16, 10, 4, 4, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 17, 0, 4, 12, -2, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 18, 6, 3, 18, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 5, 4, 2, 2, 16, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 3, 19, 17, 17, 3, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 4, 19, 16, 16, 20, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 0, 8, 3, 9, 20, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 1, 17, 2, -2, 17, 19, -2, -2, -2, -2, -2, -2, -2, -2),
                (11, 17, 7, 17, 17, 14, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 9, 4, 20, 16, 8, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 17, 2, 17, 15, 2, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 3, 3, 9, 17, 4, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 4, 0, 11, 16, 17, 15, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 17, 2, 3, 2, 16, 14, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 7, 0, 17, 5, 2, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 20, 11, 6, 3, 17, 19, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 0, 2, 17, 12, 4, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 1, 10, 2, 4, 17, 9, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 5, 16, 16, 16, 16, 5, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 4, 0, 17, 18, 17, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 5, 17, 2, 7, 0, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 12, 16, 0, 3, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 1, 1, 1, 4, 1, 19, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 18, 3, 17, 17, 1, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 17, 4, 3, 13, 18, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 3, 2, 2, 17, -2, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 1, 16, 0, 18, 3, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 20, 20, 20, 0, 10, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (20, 12, 17, 3, 4, 17, 12, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 16, 17, 0, 2, 13, 15, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 9, 4, 19, 8, 2, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 3, 1, 3, 0, 17, 6, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 20, 0, 16, 20, 14, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 3, 1, 18, 18, 1, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 15, 3, 17, 17, 17, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 0, 16, 0, 1, 1, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 16, 0, 2, 1, 20, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 15, 14, 20, 17, 15, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 6, 16, 11, 17, 17, 20, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 4, 2, 9, 1, 0, 7, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 4, 16, 17, 0, 18, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 1, 1, 1, 16, 3, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 17, 2, 17, 16, 1, 3, -2, -2, -2, -2, -2, -2, -2, -2)
                );
    constant threshold_int : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((9663676416, 988218687, 7209778183, 2994186242, 1970528513, 5856588800, 4368056838, 0, 0, 0, 0, 0, 0, 0, 0),
                (9663676416, 598020288, 7998104570, 5463109624, 6882852853, 4786012152, 1158616064, 0, 0, 0, 0, 0, 0, 0, 0),
                (1654747393, 6334658045, 11811160064, 4573687287, 4044986370, 2979571714, 9607260152, 0, 0, 0, 0, 0, 0, 0, 0),
                (9663676416, 5368709120, 5693747198, 3474510345, 1073741824, 2422798847, 11811160064, 0, 0, 0, 0, 0, 0, 0, 0),
                (2356992518, 9757571080, 3044141050, 4486000634, 12190953478, 3039430652, 5369171537654, 0, 0, 0, 0, 0, 0, 0, 0),
                (18182307851, 3766446595, 11811160064, 6723468807, 11811160064, 23341301706, 5172581371, 0, 0, 0, 0, 0, 0, 0, 0),
                (2677435647, 5082512385, 4526612405740, 23844618186, 15791554549, 3625172730, 2241661951, 0, 0, 0, 0, 0, 0, 0, 0),
                (202649664, 10641815554, 1763704831, 1073741824, 391168295422, 11811160064, 2640314889, 0, 0, 0, 0, 0, 0, 0, 0),
                (11811160064, 2659723502378, 5165178888, 9663676416, 6664748551, 2934867224848, 8047006724, 0, 0, 0, 0, 0, 0, 0, 0),
                (4267640824, 1073741824, 3348128248, 4777312761, 1073741824, 1073741824, 4161697274, 0, 0, 0, 0, 0, 0, 0, 0),
                (21076377589, 12988459004, 9663676416, 5444033032, 14312672261, 1073741824, 5024215033, 0, 0, 0, 0, 0, 0, 0, 0),
                (1073741824, 4886364665, 1073741824, 1073741824, 1073741824, 2193621239, 1073741824, 0, 0, 0, 0, 0, 0, 0, 0),
                (1212372096, 4297479165, 7763657724, 9663676416, 9663676416, 1073741824, 1073741824, 0, 0, 0, 0, 0, 0, 0, 0),
                (3339619832, 4299162105, 3572742647, 1073741824, 1073741824, 9537161218, 5745422634267, 0, 0, 0, 0, 0, 0, 0, 0),
                (2850230277, -1057912065, -606543487, 4213326840, 853608759917, 4666947004688, 11639193611, 0, 0, 0, 0, 0, 0, 0, 0),
                (11496011771, 3988871677, 230943997131, 27367833546, 5317789211804, 207186591692, 1073741824, 0, 0, 0, 0, 0, 0, 0, 0),
                (1264683136, 1073741824, 11811160064, 1058090113, 9663676416, 2182365439643, 2356954786483, 0, 0, 0, 0, 0, 0, 0, 0),
                (9286189056, 1073741824, 1073741824, 9663676416, 1073741824, 1563568112371, 4980291584, 0, 0, 0, 0, 0, 0, 0, 0),
                (875712319, 9663676416, 4588569091, 6252062581436, 4857558727026, 5368709120, 1073741824, 0, 0, 0, 0, 0, 0, 0, 0),
                (13807824905, 4246104054, 3214934011, 6059132930, 6145983374625, 615482261059, 544210124198, 0, 0, 0, 0, 0, 0, 0, 0),
                (6270847802021, 25857884106, 9663676416, 1073741824, 9663676416, 490484288, 9261023232, 0, 0, 0, 0, 0, 0, 0, 0),
                (1556086784, 1073741824, 3221225472, 1073741824, 11811160064, 1073741824, 4638900224, 0, 0, 0, 0, 0, 0, 0, 0),
                (62432223147, 5471101441, -1867847040, 9663676416, 3747389954, 1073741824, -1099700864, 0, 0, 0, 0, 0, 0, 0, 0),
                (9625927691, 9663676416, 9663676416, 3057521784196, 4170251495948, 4021077403333, 4285171506390, 0, 0, 0, 0, 0, 0, 0, 0),
                (12782760951, 477357931739, 338128503038, 7593487362, 7815891978, 3198156795, 1073741824, 0, 0, 0, 0, 0, 0, 0, 0),
                (-1092050432, 3376414473, 7649271814, 2088763521, 1073741824, 50277277794, 4852586378963, 0, 0, 0, 0, 0, 0, 0, 0),
                (4521171455, 1073741824, 5976883189, 1073741824, 1073741824, 3665269105508, 13501102070, 0, 0, 0, 0, 0, 0, 0, 0),
                (2354914806, 9663676416, 4051698179, 4959770766758, 1328204218083, 1073741824, 1073741824, 0, 0, 0, 0, 0, 0, 0, 0),
                (5230494753132, 11811160064, 9663676416, 1073741824, 6053164042, 13904117771, 4374077437, 0, 0, 0, 0, 0, 0, 0, 0),
                (1256194049, 1073741824, 6981993476, 1073741824, 1073741824, 3133145099, 1141459909784, 0, 0, 0, 0, 0, 0, 0, 0),
                (1632813057, -10336032759, 1073741824, 4655677440, 3154116608, 5775557113, 6440348149, 0, 0, 0, 0, 0, 0, 0, 0),
                (5561646589, 1073741824, 1073741824, 1073741824, 1073741824, 1073741824, 9663676416, 0, 0, 0, 0, 0, 0, 0, 0),
                (553602579872, 9663676416, 1073741824, 3854035452, 9600073727, 9663676416, 1073741824, 0, 0, 0, 0, 0, 0, 0, 0),
                (6253167762421, 3124756727, 1199389312, 1073741824, 1073741824, 9663676416, 3221225472, 0, 0, 0, 0, 0, 0, 0, 0),
                (4988755976, 30261903414, 4019419868079, 3221225472, 11811160064, 9663676416, 6347471350, 0, 0, 0, 0, 0, 0, 0, 0),
                (4674589706, 87847108650, 4821352453, 6837299721, 14315345921, 6196260498016, 1303881217, 0, 0, 0, 0, 0, 0, 0, 0),
                (5012193291, 5368709120, 1073741824, 1073741824, 3338742799490, 1073741824, 1073741824, 0, 0, 0, 0, 0, 0, 0, 0),
                (2218787063, 8361894399, 2856320777, 9663676416, 3270232766834, 1073741824, 2426183689, 0, 0, 0, 0, 0, 0, 0, 0),
                (3368733182, 2364374536, 12016680949, 9663676416, 4042703874, 160496624, 18182307851, 0, 0, 0, 0, 0, 0, 0, 0),
                (7634708482, 1073741824, 1073741824, 3373550009026, 6299845123, 9663676416, -3092323324, 0, 0, 0, 0, 0, 0, 0, 0),
                (-3358564610, 3072327675, -187030496, 4405062533456, 1493400943893, 295698431, 12387876869, 0, 0, 0, 0, 0, 0, 0, 0),
                (-4483956745, -11647794175, 613272255572, 0, 3401727335245, 5581538816, 8010930695, 0, 0, 0, 0, 0, 0, -4294967296, -4294967296),
                (8120448517, 122654474307, 9357492235, 6774793731, 1073741824, 15288238069, 9663676416, 0, 0, 0, 0, 0, 0, 0, 0),
                (3221225472, 1073741824, 4039115514, 3397385982, 10286096376, 11811160064, -753435393, 0, 0, 0, 0, 0, 0, 0, 0),
                (6141563101658, 5366961669606, 9663676416, 3552068607, 1672412033, 499734368, 5031813625, 0, 0, 0, 0, 0, 0, 0, 0),
                (4970203135, 4374572024, 9663676416, 1073741824, 9663676416, 3147578744358, -136013120, 0, 0, 0, 0, 0, 0, 0, 0),
                (3221225472, 1073741824, 4185914877, 1073741824, 2196730279887, 3221225472, 5257750530, 0, 0, 0, 0, 0, 0, 0, 0),
                (2627265275, 9663676416, 3310057465, 592607295, 1887331680675, -1625198080, 11400894458, 0, 0, 0, 0, 0, 0, 0, 0),
                (-1428524544, 1073741824, 553656641, 1073741824, 3571517958, 9663676416, 2538173887792, 0, 0, 0, 0, 0, 0, 0, 0),
                (-995301185, 1073741824, 14550787074, 2705326069, -5146292220, 4674589706, 692060160, 0, 0, 0, 0, 0, 0, 0, 0),
                (1073741824, 1073741824, 1073741824, 3374317563, 1073741824, 1073741824, 1073741824, 0, 0, 0, 0, 0, 0, 0, 0),
                (24473763894, 18308136949, 1073741824, 7996439561, 6534725632, 6276021240, 3221225472, 0, 0, 0, 0, 0, 0, 0, 0),
                (-446813696, 1073741824, -379161536, 2195718149, 9538370552, 6161452493911, 3371340398676, 0, 0, 0, 0, 0, 0, 0, 0),
                (8012735483, 890626047954, 177904205821, 9663676416, 4510037568599, 8033100285, 4937118915966, 0, 0, 0, 0, 0, 0, 0, 0),
                (6285764846210, 150994960, 4439670779, 9663676416, -1114488576, 1492504576, 4750049275, 0, 0, 0, 0, 0, 0, 0, 0),
                (2146890751, 1661148161, 1073741824, 1385922559, 3126311935, 3400622669656, 9141825542, 0, 0, 0, 0, 0, 0, 0, 0),
                (-8951519234, 4767824899, 3349151739, 0, 3353346311, 3621621586261, 5726250502, 0, 0, 0, 0, 0, 0, -4294967296, -4294967296),
                (8690332674, 1070740208796, 1073741824, 9663676416, 9663676416, 1561358106884, 3250343374582, 0, 0, 0, 0, 0, 0, 0, 0),
                (1972343551, 2132803583, 1973588735, 9663676416, 1073741824, 0, 20971524, 0, 0, 0, 0, 0, 0, -4294967296, -4294967296),
                (30639390666, 440401920, 1073741824, 5031914492, 692060160, 4580757211605, 891731050697, 0, 0, 0, 0, 0, 0, 0, 0),
                (7486832629, 1073741824, 9663676416, 3311230463, 3309145085, 2002251154247, 15288238069, 0, 0, 0, 0, 0, 0, 0, 0),
                (22460497974, 7587705863, 5368709120, 3391094779, 9468642295, 6880829430, -2637744630, 0, 0, 0, 0, 0, 0, 0, 0),
                (8012307447, 9663676416, 9663676416, 3563609119397, 1880701797359, 1073741824, 4922084361, 0, 0, 0, 0, 0, 0, 0, 0),
                (4042703874, 6616022019, 1073741824, 2636200697, 1073741824, 5368709120, 6258862073, 0, 0, 0, 0, 0, 0, 0, 0),
                (32597356520, 1021682049, 7864318980, 10145038333, 0, 7818182656, 5368709120, 0, 0, 0, 0, 0, 0, -4294967296, -4294967296),
                (1073741824, 3424648953, 1073741824, 2315255550, 5530189819, 1073741824, 9663676416, 0, 0, 0, 0, 0, 0, 0, 0),
                (2569925378, 1073741824, 11811160064, 9663676416, 2691215383708, 1073741824, 6090124297, 0, 0, 0, 0, 0, 0, 0, 0),
                (9101641720, 8529117189, 6705420281, 8514435574, 1073741824, 2883014407, 1253616909782, 0, 0, 0, 0, 0, 0, 0, 0),
                (-1487203328, -8044467711, 425994081, 1073741824, 270532607, 9663676416, 632368065, 0, 0, 0, 0, 0, 0, 0, 0),
                (5258820599, 11811160064, 6048910328, 1073741824, 1888436616847, 5144313851, 1073741824, 0, 0, 0, 0, 0, 0, 0, 0),
                (10770972672, 10468982784, 11452752903, 4042703874, 10782695420, 4198429101339, 1073741824, 0, 0, 0, 0, 0, 0, 0, 0),
                (3007876085, 1073741824, 3217971197, 6616515081, 1073741824, 2347988484, 1543125599198, 0, 0, 0, 0, 0, 0, 0, 0),
                (4571791875, 5368709120, 1073741824, 1073741824, 5513228284, 5507120647, 5368709120, 0, 0, 0, 0, 0, 0, 0, 0),
                (6055372793179, 8012735483, 7286337543, 3149922315, 1073741824, 9663676416, 1918893952, 0, 0, 0, 0, 0, 0, 0, 0),
                (562562945, -5900194, 1073741824, 10707811334, 9663676416, 3548381184, 1073741824, 0, 0, 0, 0, 0, 0, 0, 0),
                (8834549751, 1073741824, 5243754519766, 2181812978000, 1985676312811, 207186591692, 1073741824, 0, 0, 0, 0, 0, 0, 0, 0),
                (3823233020, 9663676416, 4130667510, 10798235643, 3082813451, 201326608, 4160781823, 0, 0, 0, 0, 0, 0, 0, 0),
                (2441085186, 1073741824, 2833252357, 4348998650, 1073741824, 12826451979, 4324951321687, 0, 0, 0, 0, 0, 0, 0, 0),
                (4847768070, 5173896190, 1073741824, 361333390999, 5175529480, -1312434176, 5210078218, 0, 0, 0, 0, 0, 0, 0, 0),
                (8010930695, 1302467329, 1162035713, 600409024, 9663676416, 784637568, 9663676416, 0, 0, 0, 0, 0, 0, 0, 0),
                (-10336032759, 8241807349, -7281697797, 2785017856, 4141875205, 1122141057, -5989853174, 0, 0, 0, 0, 0, 0, 0, 0),
                (9751756789, 6819938304, 9663676416, 6481002506, 1073741824, 13778288629, 14659092491, 0, 0, 0, 0, 0, 0, 0, 0),
                (121549471779, 1911519487, -13229901815, 4817112054, 6616515081, 0, -6041882623, 0, 0, 0, 0, 0, 0, -4294967296, -4294967296),
                (12270436357, 3063731963, 4383515863648, 3128694782, 2831155211, -304401151, 3435468792, 0, 0, 0, 0, 0, 0, 0, 0),
                (2007776232389, 11811160064, 11811160064, 1073741824, 10682251253, 1073741824, 1790984704, 0, 0, 0, 0, 0, 0, 0, 0),
                (1073741824, 1073741824, 9149874181, 6365383683, 9663676416, 9045016571, 1073741824, 0, 0, 0, 0, 0, 0, 0, 0),
                (8010930695, 225971503039, 6360662011, 6619608574, 7858029559, 1073741824, 1073741824, 0, 0, 0, 0, 0, 0, 0, 0),
                (2386500103, 1073741824, 11811160064, 3221225472, 1073741824, 10287626244, 10504312841, 0, 0, 0, 0, 0, 0, 0, 0),
                (4374572024, 4304202249, 1636297472, 4288758792, 8903058431, 7946108923, 1073741824, 0, 0, 0, 0, 0, 0, 0, 0),
                (4137680891, 3221225472, 4444190716, 6294604876748, 5368709120, 1073741824, -753435393, 0, 0, 0, 0, 0, 0, 0, 0),
                (297795616, 2681153285, 973599937, 14155776011, 1195376640, 934374016, 4336000704876, 0, 0, 0, 0, 0, 0, 0, 0),
                (-1750769921, 1073741824, -1736009729, 4213178363, 8587837445, 2959081220, -1735697152, 0, 0, 0, 0, 0, 0, 0, 0),
                (12162447350, 12005108740, 3891792960668, 11961960446, -52355540, 2402373636, 5057795063, 0, 0, 0, 0, 0, 0, 0, 0),
                (4919438339494, 4879105912230, 11339872250, 9671725056, 825924992, 9663676416, 13026129926, 0, 0, 0, 0, 0, 0, 0, 0),
                (6819938304, 1073741824, 1073741824, 3221225472, 5892997625, 1073741824, 1086037759, 0, 0, 0, 0, 0, 0, 0, 0),
                (2390706422, 1073741824, 3307802714083, 1073741824, 8363442691, 260046848, 11811160064, 0, 0, 0, 0, 0, 0, 0, 0),
                (5173896190, 9663676416, 2807795206, 1073741824, 2837306871, 7347539968, 1073741824, 0, 0, 0, 0, 0, 0, 0, 0),
                (173484245098, 9663676416, 224313999998, 2510290939, 6996018692, 5473566709, 14748679173, 0, 0, 0, 0, 0, 0, 0, 0),
                (1649742847, 1609037183, 1879278591, 1595972992, 4221633564099, 4140485118, 135264736, 0, 0, 0, 0, 0, 0, 0, 0),
                (828237183, 10819207173, 849957823, 6836715005, 6282449775703, -551563265, 4042703874, 0, 0, 0, 0, 0, 0, 0, 0)
                );
    constant children_left : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 13, 7, 9, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 13, 7, 9, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 13, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 13, 9, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 13, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1)
                );
    constant children_right : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 14, 8, 10, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 14, 8, 10, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 14, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 14, 10, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 14, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1)
                );
    constant value_int : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((0, 0, 0, 0, 0, 0, 0, 235596976, -1228470911, -1287112447, -1801872255, 1767209088, 1138272127, 289080288, -1357531009),
                (0, 0, 0, 0, 0, 0, 0, 993816065, -469949760, -1180154881, -469754815, 1109989503, -595058111, 113235496, -905675392),
                (0, 0, 0, 0, 0, 0, 0, 1033142656, 628609857, 120613672, -748500415, -713983552, -1118744704, 650627201, -404569695),
                (0, 0, 0, 0, 0, 0, 0, 460724511, -741477888, 773699903, -483599041, 948475201, 694625024, -252982928, 374950303),
                (0, 0, 0, 0, 0, 0, 0, 490589249, -485691264, -171469408, -703514752, -284522271, -774266049, -971990465, -538830592),
                (0, 0, 0, 0, 0, 0, 0, 145533328, 711402880, -588287744, 88561768, -699811264, -1054864704, 417164895, -881761472),
                (0, 0, 0, 0, 0, 0, 0, 528650207, -674389825, 31007080, -467707744, -629146049, -941042431, 2880274, -542738241),
                (0, 0, 0, 0, 0, 0, 0, 646137472, 214483168, -923617601, -111361680, -707007617, 283979327, 148349376, -286278208),
                (0, 0, 0, 0, 0, 0, 0, -681604481, 21836504, -97185456, 445376096, 548534465, 92579640, -194210240, -740766272),
                (0, 0, 0, 0, 0, 0, 0, -892763840, 295254881, -559530431, 630233279, 272542688, -106515848, -521839967, -848523456),
                (0, 0, 0, 0, 0, 0, 0, 106373448, -408652512, -476597985, -878455680, -518271807, -824246976, 503284833, -200810064),
                (0, 0, 0, 0, 0, 0, 0, 198648208, -1038571009, -752945344, 222117152, -713727935, -119396488, 266640800, -218032705),
                (0, 0, 0, 0, 0, 0, 0, 355108991, 648276095, -433251169, 475103615, -315002591, 10888355, -683961409, 263309312),
                (0, 0, 0, 0, 0, 0, 0, -640640960, 69798928, 383096192, 39055552, -21453464, -252335391, -726684479, 45928664),
                (0, 0, 0, 0, 0, 0, 0, 625764799, -574431488, 868215168, 192065184, 167599568, -37563556, -16279464, -218552752),
                (0, 0, 0, 0, 0, 0, 0, 49771744, -543541376, -678436927, -35255660, -1112205056, -660672449, -93818168, -455724800),
                (0, 0, 0, 0, 0, 0, 0, 72596632, 337807104, -737869248, -16009809, -270281184, -45314924, 336209632, -85536768),
                (0, 0, 0, 0, 0, 0, 0, -388681280, 36095660, -96901208, 53085916, -768483008, 704411393, 149272896, -279683200),
                (0, 0, 0, 0, 0, 0, 0, 50902332, 1028474432, 684411263, 221565152, -488166273, -30071706, -417600448, 127652344),
                (0, 0, 0, 0, 0, 0, 0, 21643584, -221545857, -590867264, 558686464, -216154097, -860556799, -1006389824, -230998047),
                (0, 0, 0, 0, 0, 0, 0, 108615776, -21208572, -494342176, -31095456, 627507201, 1554341376, -114324344, -1114355456),
                (0, 0, 0, 0, 0, 0, 0, -649963712, 559780800, -338996960, 23789468, 315894720, -124375400, -202873456, 32746798),
                (0, 0, 0, 0, 0, 0, 0, -909359935, 692307584, -1311765248, -598643520, 364657599, 72756984, 134663616, -29820724),
                (0, 0, 0, 0, 0, 0, 0, -211277968, 346351967, 114874872, -232059265, -329824031, 9568237, 174320896, -165173776),
                (0, 0, 0, 0, 0, 0, 0, 710594497, -389876288, -45473872, 56247268, -330965376, -940191616, -82128152, -338407328),
                (0, 0, 0, 0, 0, 0, 0, 242842815, 700485312, -536279201, 185150864, -992726784, -3301546, -474670880, 135306768),
                (0, 0, 0, 0, 0, 0, 0, -351534528, 59664904, 72603704, -153897504, -594021632, 71261568, -709356161, 925149313),
                (0, 0, 0, 0, 0, 0, 0, -371142272, 93877592, 790888960, 226752143, 151368928, -92983120, 133134040, -53867156),
                (0, 0, 0, 0, 0, 0, 0, -73676032, 82960720, 270855520, -9739840, 238095871, -131456824, -262827631, 167885664),
                (0, 0, 0, 0, 0, 0, 0, -46907604, -628358912, 255724320, -86817184, 166342640, -145964496, -182273168, 82217952),
                (0, 0, 0, 0, 0, 0, 0, -3393862649, 56015452, 440528864, 130273656, -11997571, -492296833, -96423056, 70775368),
                (0, 0, 0, 0, 0, 0, 0, -290040192, 215639953, -40977824, 105738368, 678435328, -400815711, -178446032, 74338344),
                (0, 0, 0, 0, 0, 0, 0, 459593376, -514605344, 653663487, -143678496, 28940856, -188266752, -592732287, -23770682),
                (0, 0, 0, 0, 0, 0, 0, 268411535, 3446383, -8758870, -254840113, 323088511, -29673956, 1157147647, 326487297),
                (0, 0, 0, 0, 0, 0, 0, 41683544, -18530672, -577333567, 554657729, -185288336, -583957953, -357404159, 94870616),
                (0, 0, 0, 0, 0, 0, 0, 124897792, -880003649, 7965247, -281944960, -764429375, 0, 237275135, -476379903),
                (0, 0, 0, 0, 0, 0, 0, 96030240, -459412927, 63627528, -50312612, -277748255, 153448560, -421478017, 31600814),
                (0, 0, 0, 0, 0, 0, 0, -141133088, 100965152, -13249586, -743485375, 614903615, 178715904, 43857552, -50346784),
                (0, 0, 0, 0, 0, 0, 0, -86189376, 188995360, -15330106, 53329944, 399835488, -133701992, -495209407, -185668160),
                (0, 0, 0, 0, 0, 0, 0, -189924992, 21230034, 3224652, 108079544, -86756904, 2240369660, 293211071, -558442559),
                (0, 0, 0, 0, 0, 0, 0, 479619969, 69090072, -443239008, 105029456, -793114560, 538400129, -4691090, 1195926271),
                (0, 0, 0, -1804297855, 0, 0, 0, -145050128, 532356639, 544122241, -78181336, -44623468, 22561352, -1804297855, -1804297855),
                (0, 0, 0, 0, 0, 0, 0, 249642560, -833950720, 16733119, -31046148, -539602047, 6129659, 405694304, -341689057),
                (0, 0, 0, 0, 0, 0, 0, 14659199, -175184464, 201762576, 775840320, -294448353, 95690168, 127319512, -8282465),
                (0, 0, 0, 0, 0, 0, 0, 7874826, -177134672, -85285096, 160670688, 136144608, 546819328, -139092704, 518928991),
                (0, 0, 0, 0, 0, 0, 0, 20994796, -38081236, -124852336, 259627728, -162531072, 57142044, -659561536, -30068206),
                (0, 0, 0, 0, 0, 0, 0, 276491936, -358626335, 103403136, -61454896, 1857678335, -116988744, -79946824, 18792348),
                (0, 0, 0, 0, 0, 0, 0, -263755505, 44564988, 524903840, 151764368, -1304889216, -336609023, 4603338, -51180456),
                (0, 0, 0, 0, 0, 0, 0, 390844384, 41797600, 10742729, -140129184, -133202824, 3335038, -86693640, 53568128),
                (0, 0, 0, 0, 0, 0, 0, 806827263, -613778177, -801286592, 895103745, -5607, -385218784, 515861665, -347602623),
                (0, 0, 0, 0, 0, 0, 0, 273070881, -12525788, -799796928, -133746424, -581014719, 262712352, 169932528, -48270604),
                (0, 0, 0, 0, 0, 0, 0, 6266131, -47544272, 3836913, 285129120, -81785816, 486272160, 317367329, -268426095),
                (0, 0, 0, 0, 0, 0, 0, -236933679, 31689612, 171207168, -91885784, -117832528, -846422208, -31670376, 13553876),
                (0, 0, 0, 0, 0, 0, 0, -373596032, 444895360, -93910944, 15050565, 882639296, -615013055, 39078540, -66244100),
                (0, 0, 0, 0, 0, 0, 0, -345583233, 24422312, 111580568, 905307, 1125574911, 290984831, -945029441, 30639732),
                (0, 0, 0, 0, 0, 0, 0, 2081440, -113018240, 184938896, -63982072, -113983824, 62227048, -429741888, 62933260),
                (0, 0, 0, 0, 0, 0, 0, 0, -1815509760, 63452132, -30494944, -75231472, 6792280, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, -319975648, 374884992, 57617896, -28782290, -114851840, 42442388, -69488088, -408384255),
                (0, 0, 0, 0, 0, -2115489919, 0, -303231071, 357840129, 397062176, -17784232, 244879680, -3740538, -2115489919, -2115489919),
                (0, 0, 0, 0, 0, 0, 0, -40747424, -346449921, 92765736, -291427, -158288880, 1036388225, 851803521, -486437057),
                (0, 0, 0, 0, 0, 0, 0, -248127184, 131966496, 104922424, -13283540, -229211152, -23608068, -28297086, 154084272),
                (0, 0, 0, 0, 0, 0, 0, 20923756, -7683337, -256467296, 136376528, -216688528, 598291264, -598993920, 126267856),
                (0, 0, 0, 0, 0, 0, 0, -164461088, 122259664, 215592721, -84519424, -243328016, 14841220, 234286272, -273874433),
                (0, 0, 0, 0, 0, 0, 0, -17601976, 97709456, 7117192, -99965672, 37790164, -267342097, -1384222, 244413633),
                (0, 0, 0, 0, 0, 0, 0, -1278364288, -157447184, 4441241, 572471937, 427121952, -48808892, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, -12267895, 67692328, -346101631, 15719729, -142709872, 37857984, 179767856, 18677944),
                (0, 0, 0, 0, 0, 0, 0, 34158744, 407903616, 66278612, -107714224, -105340240, 36523816, 214450032, -23692902),
                (0, 0, 0, 0, 0, 0, 0, -1489413, 528812288, 144502896, -296442111, 151690672, -164984112, -334878624, 144358832),
                (0, 0, 0, 0, 0, 0, 0, 130412336, -1173622528, -306507393, 847683329, 32131164, -119646928, 135704512, 355090),
                (0, 0, 0, 0, 0, 0, 0, -19837464, -266843825, 395472703, 39730280, 55565848, 279278208, 16458912, -44078332),
                (0, 0, 0, 0, 0, 0, 0, -7099181, 39383276, -71932776, -494987553, 344418111, 0, 240357760, -519920192),
                (0, 0, 0, 0, 0, 0, 0, 375303904, -91577816, -421319775, 48796536, -58546976, -540953345, -39308200, 3537425),
                (0, 0, 0, 0, 0, 0, 0, 755909951, -213786768, 6808059, -120831248, -326718401, 15960787, 297213023, 7191838),
                (0, 0, 0, 0, 0, 0, 0, 15398218, -60800524, -28610406, 51995948, 223244527, 32728872, -824101888, -35563480),
                (0, 0, 0, 0, 0, 0, 0, -9333913, 85510720, -169764256, -5674410, 102141416, 2925670, -329700736, 12390364),
                (0, 0, 0, 0, 0, 0, 0, -387507935, 165650144, 105580136, -22628184, -399196607, 1488489, -373249952, -57537928),
                (0, 0, 0, 0, 0, 0, 0, -92384336, 567583424, -33590780, 195290480, -909381056, -134795536, 392250273, -3368223),
                (0, 0, 0, 0, 0, 0, 0, -244525983, 383953760, -272766080, -19931392, 156411744, -369230272, -25217326, 36124132),
                (0, 0, 0, 0, 0, 0, 0, 555012225, 11745553, -1639794432, -6581118, 0, -613210880, -330267712, 337173569),
                (0, 0, 0, 0, 0, 0, 0, -16126404, 98716912, 12530130, -192271456, 3549026, -104219000, 44974400, 321164224),
                (0, 0, 0, 0, 0, 0, 0, 400004448, -1322876543, -197925472, 1167571456, 151599600, 688913856, -302048128, -1606621),
                (0, 0, 0, 0, 0, 0, 0, 24171510, -237183249, -283756128, -3913269, 16126165, -104391144, -27418642, 75781424),
                (0, 0, 0, 0, 0, -1348171903, 0, 8152381, -867143873, -158772304, 861385984, 277676289, 973828, -1348171903, -1348171903),
                (0, 0, 0, 0, 0, 0, 0, 61672084, -2064495, 125424232, -94986488, -987177664, 301133727, 1337290881, 0),
                (0, 0, 0, 0, 0, 0, 0, 296832287, -72728792, 265392208, -40497228, 8647040, 104202968, -251563968, -28707098),
                (0, 0, 0, 0, 0, 0, 0, 655760192, 4191193348, -229759855, 83487912, 1825479, -254794000, -522074080, 105269080),
                (0, 0, 0, 0, 0, 0, 0, 491874719, -234890479, -9350645, -309636225, 37510988, -108094136, 193799136, -38181644),
                (0, 0, 0, 0, 0, 0, 0, 132097256, 7905757, 142572224, -47657912, -60571964, 47108300, 53653364, -89363088),
                (0, 0, 0, 0, 0, 0, 0, -3618963, 441464929, -313213823, -33170690, 139968352, -64687904, 62497732, -165886720),
                (0, 0, 0, 0, 0, 0, 0, 1597598848, -764912703, -212031440, -4656902, -272381120, 15120582, 137788880, 7848939),
                (0, 0, 0, 0, 0, 0, 0, -102668672, -421845183, -336712319, 62136604, -3920901, -231348416, -19131638, 73329696),
                (0, 0, 0, 0, 0, 0, 0, -100461224, 144169280, -615024321, 100339960, -99068280, 1147537151, -1921939584, 5669168),
                (0, 0, 0, 0, 0, 0, 0, 1209168, 231536097, 64117296, -286952256, 106903040, -165665920, -351901984, 520489567),
                (0, 0, 0, 0, 0, 0, 0, -14176496, 23671002, 320139872, 2555311, 13162557, -101931616, -348342848, 262456544),
                (0, 0, 0, 0, 0, 0, 0, 188065760, -3942534, 390358911, 20098498, 295579647, -240070240, -200374080, -25954724),
                (0, 0, 0, 0, 0, 0, 0, -194010528, -7576310, 29619752, -443905153, 106532312, -56571900, 27732944, -62080392),
                (0, 0, 0, 0, 0, 0, 0, -125813584, 70925048, 56805396, 577532864, -345841023, 179677712, -26484630, 14630228),
                (0, 0, 0, 0, 0, 0, 0, -882444032, 0, 648135104, -294779039, -44587200, 468527713, -308286, -221781185),
                (0, 0, 0, 0, 0, 0, 0, -2861942, 379271425, -367178464, -42106244, 181574496, -123286968, -203001536, 9053432),
                (0, 0, 0, 0, 0, 0, 0, 66955488, -181575376, 637482368, -2000368640, -1501705600, 71109400, -11161875, 16761999)
                );
    constant parent : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 4, 4, 5, 5, 6, 6, 3, 3),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 4, 4, 5, 5, 6, 6, 3, 3),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 6, 6, 5, 5),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 5, 5, 6, 6, 4, 4),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 6, 6, 5, 5),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6)
                );
    constant depth : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3)
                );
    constant iLeaf : intArray2D(nTrees-1 downto 0)(nLeaves-1 downto 0) := ((7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14)
                );
    constant value : tyArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := to_tyArray2D(value_int);
      constant threshold : txArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := to_txArray2D(threshold_int);
end Arrays0;