library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_misc.all;
  use ieee.numeric_std.all;

  use work.Constants.all;
  use work.Types.all;
  package Arrays0 is

    constant initPredict : ty := to_ty(0);
    constant feature : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((4, 1, 0, 3, 1, 0, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 1, 0, 0, 17, 3, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 4, 0, 3, 3, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 19, 0, 0, 15, 2, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 1, 3, 0, 3, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 3, 4, 17, 4, 18, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 16, 18, 18, 1, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 17, 5, 16, 4, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 16, 3, 4, 17, 16, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 7, 1, 17, 6, 5, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 0, 4, 3, 2, 5, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (7, 17, 6, 5, 12, 17, 13, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 3, 17, 20, 20, 7, 13, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 17, 1, 7, 14, 0, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 2, 1, 1, 16, 16, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 1, 16, 18, 16, 16, 10, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 10, 4, 1, 4, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 6, 14, 4, 7, 16, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 20, 17, 16, 16, 20, 12, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 1, 17, 3, 16, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 18, 4, 5, 4, 1, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 5, 19, 9, 4, 10, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 2, 1, 4, 3, 5, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 4, 4, 16, 16, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 16, 16, 0, 2, 17, 10, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 17, 3, 17, 13, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 7, 18, 13, 13, 16, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 4, 17, 16, 16, 5, 14, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 4, 4, 8, 2, 18, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 8, 2, 10, 5, 17, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 3, 12, 18, 17, 17, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 7, 14, 10, 11, 15, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 4, 10, 0, 2, 20, 8, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 17, 1, 5, 9, 4, 19, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 18, 16, 19, 4, 19, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 16, 17, 0, 2, 16, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 20, 15, 13, 16, 12, 13, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 2, 17, 4, 16, 5, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 2, 18, 4, 3, 3, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 6, 6, 16, 17, 20, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 17, 0, 16, 16, 17, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 2, 16, -2, 16, 2, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 16, 17, 2, 10, 18, 19, -2, -2, -2, -2, -2, -2, -2, -2),
                (19, 11, 17, 17, 2, 4, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 16, 4, 1, 1, 1, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 3, 19, 9, 4, 16, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (19, 9, 17, 10, 16, 20, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 4, 0, 1, 16, 1, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 13, 1, 5, 3, 4, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 6, 2, 18, 0, 1, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (8, 10, 5, 17, 5, 9, 9, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 18, 6, 17, 17, 0, 20, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 10, 1, 17, 0, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 16, 16, 4, 16, 2, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 17, 17, 4, 2, 2, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 1, 15, 1, 3, 16, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 17, -2, 17, 16, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 16, 10, 4, 4, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 17, 0, 4, 12, -2, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 18, 6, 3, 18, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 5, 4, 2, 2, 16, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 3, 19, 17, 17, 3, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 4, 19, 16, 16, 20, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 0, 8, 3, 9, 20, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 1, 17, 2, -2, 17, 19, -2, -2, -2, -2, -2, -2, -2, -2),
                (11, 17, 7, 17, 17, 14, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 9, 4, 20, 16, 8, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 17, 2, 17, 15, 2, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 3, 3, 9, 17, 4, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 4, 0, 11, 16, 17, 15, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 17, 2, 3, 2, 16, 14, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 7, 0, 17, 5, 2, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 20, 11, 6, 3, 17, 19, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 0, 2, 17, 12, 4, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 1, 10, 2, 4, 17, 9, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 5, 16, 16, 16, 16, 5, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 4, 0, 17, 18, 17, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 5, 17, 2, 7, 0, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 12, 16, 0, 3, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 1, 1, 1, 4, 1, 19, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 18, 3, 17, 17, 1, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 17, 4, 3, 13, 18, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 3, 2, 2, 17, -2, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 1, 16, 0, 18, 3, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 20, 20, 20, 0, 10, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (20, 12, 17, 3, 4, 17, 12, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 16, 17, 0, 2, 13, 15, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 9, 4, 19, 8, 2, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 3, 1, 3, 0, 17, 6, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 20, 0, 16, 20, 14, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 3, 1, 18, 18, 1, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 15, 3, 17, 17, 17, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 0, 16, 0, 1, 1, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 16, 0, 2, 1, 20, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 15, 14, 20, 17, 15, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 6, 16, 11, 17, 17, 20, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 4, 2, 9, 1, 0, 7, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 4, 16, 17, 0, 18, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 1, 1, 1, 16, 3, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 17, 2, 17, 16, 1, 3, -2, -2, -2, -2, -2, -2, -2, -2)
                );
    constant threshold_int : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((294912, 30158, 220025, 91375, 60136, 178729, 133303, 0, 0, 0, 0, 0, 0, 0, 0),
                (294912, 18250, 244083, 166721, 210048, 146057, 35358, 0, 0, 0, 0, 0, 0, 0, 0),
                (50499, 193318, 360448, 139578, 123443, 90929, 293190, 0, 0, 0, 0, 0, 0, 0, 0),
                (294912, 163840, 173759, 106034, 32768, 73938, 360448, 0, 0, 0, 0, 0, 0, 0, 0),
                (71930, 297777, 92900, 136902, 372038, 92756, 163854112, 0, 0, 0, 0, 0, 0, 0, 0),
                (554880, 114943, 360448, 205184, 360448, 712320, 157855, 0, 0, 0, 0, 0, 0, 0, 0),
                (81709, 155106, 138141248, 727680, 481920, 110631, 68410, 0, 0, 0, 0, 0, 0, 0, 0),
                (6184, 324762, 53824, 32768, 11937509, 360448, 80576, 0, 0, 0, 0, 0, 0, 0, 0),
                (360448, 81168320, 157629, 294912, 203392, 89565040, 245575, 0, 0, 0, 0, 0, 0, 0, 0),
                (130238, 32768, 102177, 145792, 32768, 32768, 127005, 0, 0, 0, 0, 0, 0, 0, 0),
                (643200, 396376, 294912, 166139, 436788, 32768, 153327, 0, 0, 0, 0, 0, 0, 0, 0),
                (32768, 149120, 32768, 32768, 32768, 66944, 32768, 0, 0, 0, 0, 0, 0, 0, 0),
                (36999, 131149, 236928, 294912, 294912, 32768, 32768, 0, 0, 0, 0, 0, 0, 0, 0),
                (101917, 131200, 109031, 32768, 32768, 291051, 175336384, 0, 0, 0, 0, 0, 0, 0, 0),
                (86982, -32285, -18510, 128581, 26050072, 142423920, 355200, 0, 0, 0, 0, 0, 0, 0, 0),
                (350830, 121731, 7047851, 835200, 162286048, 6322833, 32768, 0, 0, 0, 0, 0, 0, 0, 0),
                (38595, 32768, 360448, 32290, 294912, 66600508, 71928552, 0, 0, 0, 0, 0, 0, 0, 0),
                (283392, 32768, 32768, 294912, 32768, 47716312, 151986, 0, 0, 0, 0, 0, 0, 0, 0),
                (26725, 294912, 140032, 190797808, 148240928, 163840, 32768, 0, 0, 0, 0, 0, 0, 0, 0),
                (421381, 129581, 98112, 184910, 187560528, 18783028, 16607975, 0, 0, 0, 0, 0, 0, 0, 0),
                (191371088, 789120, 294912, 32768, 294912, 14968, 282624, 0, 0, 0, 0, 0, 0, 0, 0),
                (47488, 32768, 98304, 32768, 360448, 32768, 141568, 0, 0, 0, 0, 0, 0, 0, 0),
                (1905280, 166965, -57002, 294912, 114361, 32768, -33560, 0, 0, 0, 0, 0, 0, 0, 0),
                (293760, 294912, 294912, 93308160, 127265976, 122713544, 130773056, 0, 0, 0, 0, 0, 0, 0, 0),
                (390099, 14567808, 10318863, 231735, 238522, 97600, 32768, 0, 0, 0, 0, 0, 0, 0, 0),
                (-33327, 103040, 233437, 63744, 32768, 1534341, 148089184, 0, 0, 0, 0, 0, 0, 0, 0),
                (137975, 32768, 182400, 32768, 32768, 111855136, 412021, 0, 0, 0, 0, 0, 0, 0, 0),
                (71866, 294912, 123648, 151360192, 40533576, 32768, 32768, 0, 0, 0, 0, 0, 0, 0, 0),
                (159622032, 360448, 294912, 32768, 184728, 424320, 133486, 0, 0, 0, 0, 0, 0, 0, 0),
                (38336, 32768, 213074, 32768, 32768, 95616, 34834592, 0, 0, 0, 0, 0, 0, 0, 0),
                (49830, -315431, 32768, 142080, 96256, 176256, 196544, 0, 0, 0, 0, 0, 0, 0, 0),
                (169728, 32768, 32768, 32768, 32768, 32768, 294912, 0, 0, 0, 0, 0, 0, 0, 0),
                (16894610, 294912, 32768, 117616, 292971, 294912, 32768, 0, 0, 0, 0, 0, 0, 0, 0),
                (190831536, 95360, 36602, 32768, 32768, 294912, 98304, 0, 0, 0, 0, 0, 0, 0, 0),
                (152245, 923520, 122662960, 98304, 360448, 294912, 193709, 0, 0, 0, 0, 0, 0, 0, 0),
                (142657, 2680881, 147136, 208658, 436870, 189094864, 39791, 0, 0, 0, 0, 0, 0, 0, 0),
                (152960, 163840, 32768, 32768, 101890344, 32768, 32768, 0, 0, 0, 0, 0, 0, 0, 0),
                (67712, 255185, 87168, 294912, 99799584, 32768, 74041, 0, 0, 0, 0, 0, 0, 0, 0),
                (102806, 72155, 366720, 294912, 123374, 4898, 554880, 0, 0, 0, 0, 0, 0, 0, 0),
                (232993, 32768, 32768, 102952576, 192256, 294912, -94370, 0, 0, 0, 0, 0, 0, 0, 0),
                (-102495, 93760, -5708, 134431840, 45574980, 9024, 378048, 0, 0, 0, 0, 0, 0, 0, 0),
                (-136840, -355462, 18715584, 0, 103812480, 170335, 244474, 0, 0, 0, 0, 0, 0, -131072, -131072),
                (247816, 3743118, 285568, 206750, 32768, 466560, 294912, 0, 0, 0, 0, 0, 0, 0, 0),
                (98304, 32768, 123264, 103680, 313907, 360448, -22993, 0, 0, 0, 0, 0, 0, 0, 0),
                (187425632, 163786672, 294912, 108401, 51038, 15251, 153559, 0, 0, 0, 0, 0, 0, 0, 0),
                (151679, 133501, 294912, 32768, 294912, 96056480, -4151, 0, 0, 0, 0, 0, 0, 0, 0),
                (98304, 32768, 127744, 32768, 67038888, 98304, 160454, 0, 0, 0, 0, 0, 0, 0, 0),
                (80178, 294912, 101015, 18085, 57596792, -49597, 347928, 0, 0, 0, 0, 0, 0, 0, 0),
                (-43595, 32768, 16896, 32768, 108994, 294912, 77458920, 0, 0, 0, 0, 0, 0, 0, 0),
                (-30374, 32768, 444055, 82560, -157052, 142657, 21120, 0, 0, 0, 0, 0, 0, 0, 0),
                (32768, 32768, 32768, 102976, 32768, 32768, 32768, 0, 0, 0, 0, 0, 0, 0, 0),
                (746880, 558720, 32768, 244032, 199424, 191529, 98304, 0, 0, 0, 0, 0, 0, 0, 0),
                (-13636, 32768, -11571, 67008, 291088, 188032608, 102885144, 0, 0, 0, 0, 0, 0, 0, 0),
                (244529, 27179750, 5429205, 294912, 137635424, 245151, 150668912, 0, 0, 0, 0, 0, 0, 0, 0),
                (191826320, 4608, 135488, 294912, -34011, 45548, 144960, 0, 0, 0, 0, 0, 0, 0, 0),
                (65518, 50694, 32768, 42295, 95407, 103778768, 278986, 0, 0, 0, 0, 0, 0, 0, 0),
                (-273179, 145502, 102208, 0, 102336, 110523120, 174751, 0, 0, 0, 0, 0, 0, -131072, -131072),
                (265208, 32676398, 32768, 294912, 294912, 47648868, 99192608, 0, 0, 0, 0, 0, 0, 0, 0),
                (60191, 65088, 60229, 294912, 32768, 0, 640, 0, 0, 0, 0, 0, 0, -131072, -131072),
                (935040, 13440, 32768, 153562, 21120, 139793616, 27213472, 0, 0, 0, 0, 0, 0, 0, 0),
                (228480, 32768, 294912, 101051, 100987, 61103856, 466560, 0, 0, 0, 0, 0, 0, 0, 0),
                (685440, 231558, 163840, 103488, 288960, 209986, -80498, 0, 0, 0, 0, 0, 0, 0, 0),
                (244516, 294912, 294912, 108752720, 57394464, 32768, 150210, 0, 0, 0, 0, 0, 0, 0, 0),
                (123374, 201905, 32768, 80450, 32768, 163840, 191005, 0, 0, 0, 0, 0, 0, 0, 0),
                (994792, 31179, 240000, 309602, 0, 238592, 163840, 0, 0, 0, 0, 0, 0, -131072, -131072),
                (32768, 104512, 32768, 70656, 168768, 32768, 294912, 0, 0, 0, 0, 0, 0, 0, 0),
                (78428, 32768, 360448, 294912, 82129376, 32768, 185856, 0, 0, 0, 0, 0, 0, 0, 0),
                (277760, 260288, 204633, 259840, 32768, 87983, 38257352, 0, 0, 0, 0, 0, 0, 0, 0),
                (-45386, -245498, 13000, 32768, 8256, 294912, 19298, 0, 0, 0, 0, 0, 0, 0, 0),
                (160486, 360448, 184598, 32768, 57630512, 156992, 32768, 0, 0, 0, 0, 0, 0, 0, 0),
                (328704, 319488, 349510, 123374, 329062, 128125888, 32768, 0, 0, 0, 0, 0, 0, 0, 0),
                (91793, 32768, 98205, 201920, 32768, 71655, 47092456, 0, 0, 0, 0, 0, 0, 0, 0),
                (139520, 163840, 32768, 32768, 168250, 168064, 163840, 0, 0, 0, 0, 0, 0, 0, 0),
                (184795312, 244529, 222361, 96128, 32768, 294912, 58560, 0, 0, 0, 0, 0, 0, 0, 0),
                (17168, -180, 32768, 326776, 294912, 108288, 32768, 0, 0, 0, 0, 0, 0, 0, 0),
                (269609, 32768, 160026688, 66583648, 60598032, 6322833, 32768, 0, 0, 0, 0, 0, 0, 0, 0),
                (116676, 294912, 126058, 329536, 94080, 6144, 126977, 0, 0, 0, 0, 0, 0, 0, 0),
                (74496, 32768, 86464, 132721, 32768, 391432, 131987040, 0, 0, 0, 0, 0, 0, 0, 0),
                (147942, 157895, 32768, 11027020, 157945, -40052, 158999, 0, 0, 0, 0, 0, 0, 0, 0),
                (244474, 39748, 35463, 18323, 294912, 23945, 294912, 0, 0, 0, 0, 0, 0, 0, 0),
                (-315431, 251520, -222220, 84992, 126400, 34245, -182796, 0, 0, 0, 0, 0, 0, 0, 0),
                (297600, 208128, 294912, 197785, 32768, 420480, 447360, 0, 0, 0, 0, 0, 0, 0, 0),
                (3709396, 58335, -403745, 147007, 201920, 0, -184384, 0, 0, 0, 0, 0, 0, -131072, -131072),
                (374464, 93498, 133774288, 95480, 86400, -9290, 104842, 0, 0, 0, 0, 0, 0, 0, 0),
                (61272468, 360448, 360448, 32768, 325996, 32768, 54657, 0, 0, 0, 0, 0, 0, 0, 0),
                (32768, 32768, 279232, 194256, 294912, 276032, 32768, 0, 0, 0, 0, 0, 0, 0, 0),
                (244474, 6896103, 194112, 202014, 239808, 32768, 32768, 0, 0, 0, 0, 0, 0, 0, 0),
                (72830, 32768, 360448, 98304, 32768, 313953, 320566, 0, 0, 0, 0, 0, 0, 0, 0),
                (133501, 131354, 49936, 130883, 271700, 242496, 32768, 0, 0, 0, 0, 0, 0, 0, 0),
                (126272, 98304, 135626, 192096096, 163840, 32768, -22993, 0, 0, 0, 0, 0, 0, 0, 0),
                (9088, 81822, 29712, 432000, 36480, 28515, 132324240, 0, 0, 0, 0, 0, 0, 0, 0),
                (-53429, 32768, -52979, 128576, 262080, 90304, -52969, 0, 0, 0, 0, 0, 0, 0, 0),
                (371168, 366367, 118768096, 365050, -1598, 73315, 154352, 0, 0, 0, 0, 0, 0, 0, 0),
                (150129344, 148898496, 346065, 295158, 25205, 294912, 397526, 0, 0, 0, 0, 0, 0, 0, 0),
                (208128, 32768, 32768, 98304, 179840, 32768, 33143, 0, 0, 0, 0, 0, 0, 0, 0),
                (72959, 32768, 100946128, 32768, 255232, 7936, 360448, 0, 0, 0, 0, 0, 0, 0, 0),
                (157895, 294912, 85687, 32768, 86588, 224229, 32768, 0, 0, 0, 0, 0, 0, 0, 0),
                (5294319, 294912, 6845520, 76608, 213502, 167040, 450094, 0, 0, 0, 0, 0, 0, 0, 0),
                (50346, 49104, 57351, 48705, 128834032, 126358, 4128, 0, 0, 0, 0, 0, 0, 0, 0),
                (25276, 330176, 25939, 208640, 191725152, -16832, 123374, 0, 0, 0, 0, 0, 0, 0, 0)
                );
    constant children_left : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 13, 7, 9, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 13, 7, 9, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 13, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 13, 9, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 13, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1)
                );
    constant children_right : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 14, 8, 10, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 14, 8, 10, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 14, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 14, 10, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 14, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1)
                );
    constant value_int : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((0, 0, 0, 0, 0, 0, 0, 7190, -37490, -39280, -54989, 53931, 34737, 8822, -41429),
                (0, 0, 0, 0, 0, 0, 0, 30329, -14342, -36015, -14336, 33874, -18160, 3456, -27639),
                (0, 0, 0, 0, 0, 0, 0, 31529, 19184, 3681, -22842, -21789, -34141, 19856, -12346),
                (0, 0, 0, 0, 0, 0, 0, 14060, -22628, 23611, -14758, 28945, 21198, -7720, 11443),
                (0, 0, 0, 0, 0, 0, 0, 14972, -14822, -5233, -21470, -8683, -23629, -29663, -16444),
                (0, 0, 0, 0, 0, 0, 0, 4441, 21710, -17953, 2703, -21357, -32192, 12731, -26909),
                (0, 0, 0, 0, 0, 0, 0, 16133, -20581, 946, -14273, -19200, -28718, 88, -16563),
                (0, 0, 0, 0, 0, 0, 0, 19719, 6546, -28187, -3398, -21576, 8666, 4527, -8737),
                (0, 0, 0, 0, 0, 0, 0, -20801, 666, -2966, 13592, 16740, 2825, -5927, -22606),
                (0, 0, 0, 0, 0, 0, 0, -27245, 9010, -17076, 19233, 8317, -3251, -15925, -25895),
                (0, 0, 0, 0, 0, 0, 0, 3246, -12471, -14545, -26808, -15816, -25154, 15359, -6128),
                (0, 0, 0, 0, 0, 0, 0, 6062, -31695, -22978, 6778, -21781, -3644, 8137, -6654),
                (0, 0, 0, 0, 0, 0, 0, 10837, 19784, -13222, 14499, -9613, 332, -20873, 8036),
                (0, 0, 0, 0, 0, 0, 0, -19551, 2130, 11691, 1192, -655, -7701, -22177, 1402),
                (0, 0, 0, 0, 0, 0, 0, 19097, -17530, 26496, 5861, 5115, -1146, -497, -6670),
                (0, 0, 0, 0, 0, 0, 0, 1519, -16588, -20704, -1076, -33942, -20162, -2863, -13908),
                (0, 0, 0, 0, 0, 0, 0, 2215, 10309, -22518, -489, -8248, -1383, 10260, -2610),
                (0, 0, 0, 0, 0, 0, 0, -11862, 1102, -2957, 1620, -23452, 21497, 4555, -8535),
                (0, 0, 0, 0, 0, 0, 0, 1553, 31387, 20887, 6762, -14898, -918, -12744, 3896),
                (0, 0, 0, 0, 0, 0, 0, 661, -6761, -18032, 17050, -6596, -26262, -30713, -7050),
                (0, 0, 0, 0, 0, 0, 0, 3315, -647, -15086, -949, 19150, 47435, -3489, -34007),
                (0, 0, 0, 0, 0, 0, 0, -19835, 17083, -10345, 726, 9640, -3796, -6191, 999),
                (0, 0, 0, 0, 0, 0, 0, -27751, 21128, -40032, -18269, 11128, 2220, 4110, -910),
                (0, 0, 0, 0, 0, 0, 0, -6448, 10570, 3506, -7082, -10065, 292, 5320, -5041),
                (0, 0, 0, 0, 0, 0, 0, 21686, -11898, -1388, 1717, -10100, -28692, -2506, -10327),
                (0, 0, 0, 0, 0, 0, 0, 7411, 21377, -16366, 5650, -30296, -101, -14486, 4129),
                (0, 0, 0, 0, 0, 0, 0, -10728, 1821, 2216, -4697, -18128, 2175, -21648, 28233),
                (0, 0, 0, 0, 0, 0, 0, -11326, 2865, 24136, 6920, 4619, -2838, 4063, -1644),
                (0, 0, 0, 0, 0, 0, 0, -2248, 2532, 8266, -297, 7266, -4012, -8021, 5123),
                (0, 0, 0, 0, 0, 0, 0, -1432, -19176, 7804, -2649, 5076, -4454, -5563, 2509),
                (0, 0, 0, 0, 0, 0, 0, -103572, 1709, 13444, 3976, -366, -15024, -2943, 2160),
                (0, 0, 0, 0, 0, 0, 0, -8851, 6581, -1251, 3227, 20704, -12232, -5446, 2269),
                (0, 0, 0, 0, 0, 0, 0, 14026, -15705, 19948, -4385, 883, -5745, -18089, -725),
                (0, 0, 0, 0, 0, 0, 0, 8191, 105, -267, -7777, 9860, -906, 35313, 9964),
                (0, 0, 0, 0, 0, 0, 0, 1272, -566, -17619, 16927, -5655, -17821, -10907, 2895),
                (0, 0, 0, 0, 0, 0, 0, 3812, -26856, 243, -8604, -23329, 0, 7241, -14538),
                (0, 0, 0, 0, 0, 0, 0, 2931, -14020, 1942, -1535, -8476, 4683, -12862, 964),
                (0, 0, 0, 0, 0, 0, 0, -4307, 3081, -404, -22689, 18765, 5454, 1338, -1536),
                (0, 0, 0, 0, 0, 0, 0, -2630, 5768, -468, 1628, 12202, -4080, -15113, -5666),
                (0, 0, 0, 0, 0, 0, 0, -5796, 648, 98, 3298, -2648, 68371, 8948, -17042),
                (0, 0, 0, 0, 0, 0, 0, 14637, 2108, -13527, 3205, -24204, 16431, -143, 36497),
                (0, 0, 0, -55063, 0, 0, 0, -4427, 16246, 16605, -2386, -1362, 689, -55063, -55063),
                (0, 0, 0, 0, 0, 0, 0, 7618, -25450, 511, -947, -16467, 187, 12381, -10428),
                (0, 0, 0, 0, 0, 0, 0, 447, -5346, 6157, 23677, -8986, 2920, 3885, -253),
                (0, 0, 0, 0, 0, 0, 0, 240, -5406, -2603, 4903, 4155, 16688, -4245, 15836),
                (0, 0, 0, 0, 0, 0, 0, 641, -1162, -3810, 7923, -4960, 1744, -20128, -918),
                (0, 0, 0, 0, 0, 0, 0, 8438, -10944, 3156, -1875, 56692, -3570, -2440, 573),
                (0, 0, 0, 0, 0, 0, 0, -8049, 1360, 16019, 4631, -39822, -10272, 140, -1562),
                (0, 0, 0, 0, 0, 0, 0, 11928, 1276, 328, -4276, -4065, 102, -2646, 1635),
                (0, 0, 0, 0, 0, 0, 0, 24622, -18731, -24453, 27316, 0, -11756, 15743, -10608),
                (0, 0, 0, 0, 0, 0, 0, 8333, -382, -24408, -4082, -17731, 8017, 5186, -1473),
                (0, 0, 0, 0, 0, 0, 0, 191, -1451, 117, 8701, -2496, 14840, 9685, -8192),
                (0, 0, 0, 0, 0, 0, 0, -7231, 967, 5225, -2804, -3596, -25831, -967, 414),
                (0, 0, 0, 0, 0, 0, 0, -11401, 13577, -2866, 459, 26936, -18769, 1193, -2022),
                (0, 0, 0, 0, 0, 0, 0, -10546, 745, 3405, 28, 34350, 8880, -28840, 935),
                (0, 0, 0, 0, 0, 0, 0, 64, -3449, 5644, -1953, -3479, 1899, -13115, 1921),
                (0, 0, 0, 0, 0, 0, 0, 0, -55405, 1936, -931, -2296, 207, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, -9765, 11441, 1758, -878, -3505, 1295, -2121, -12463),
                (0, 0, 0, 0, 0, -64560, 0, -9254, 10920, 12117, -543, 7473, -114, -64560, -64560),
                (0, 0, 0, 0, 0, 0, 0, -1244, -10573, 2831, -9, -4831, 31628, 25995, -14845),
                (0, 0, 0, 0, 0, 0, 0, -7572, 4027, 3202, -405, -6995, -720, -864, 4702),
                (0, 0, 0, 0, 0, 0, 0, 639, -234, -7827, 4162, -6613, 18258, -18280, 3853),
                (0, 0, 0, 0, 0, 0, 0, -5019, 3731, 6579, -2579, -7426, 453, 7150, -8358),
                (0, 0, 0, 0, 0, 0, 0, -537, 2982, 217, -3051, 1153, -8159, -42, 7459),
                (0, 0, 0, 0, 0, 0, 0, -39013, -4805, 136, 17470, 13035, -1490, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, -374, 2066, -10562, 480, -4355, 1155, 5486, 570),
                (0, 0, 0, 0, 0, 0, 0, 1042, 12448, 2023, -3287, -3215, 1115, 6544, -723),
                (0, 0, 0, 0, 0, 0, 0, -45, 16138, 4410, -9047, 4629, -5035, -10220, 4405),
                (0, 0, 0, 0, 0, 0, 0, 3980, -35816, -9354, 25869, 981, -3651, 4141, 11),
                (0, 0, 0, 0, 0, 0, 0, -605, -8143, 12069, 1212, 1696, 8523, 502, -1345),
                (0, 0, 0, 0, 0, 0, 0, -217, 1202, -2195, -15106, 10511, 0, 7335, -15867),
                (0, 0, 0, 0, 0, 0, 0, 11453, -2795, -12858, 1489, -1787, -16509, -1200, 108),
                (0, 0, 0, 0, 0, 0, 0, 23069, -6524, 208, -3687, -9971, 487, 9070, 219),
                (0, 0, 0, 0, 0, 0, 0, 470, -1855, -873, 1587, 6813, 999, -25150, -1085),
                (0, 0, 0, 0, 0, 0, 0, -285, 2610, -5181, -173, 3117, 89, -10062, 378),
                (0, 0, 0, 0, 0, 0, 0, -11826, 5055, 3222, -691, -12183, 45, -11391, -1756),
                (0, 0, 0, 0, 0, 0, 0, -2819, 17321, -1025, 5960, -27752, -4114, 11971, -103),
                (0, 0, 0, 0, 0, 0, 0, -7462, 11717, -8324, -608, 4773, -11268, -770, 1102),
                (0, 0, 0, 0, 0, 0, 0, 16938, 358, -50043, -201, 0, -18714, -10079, 10290),
                (0, 0, 0, 0, 0, 0, 0, -492, 3013, 382, -5868, 108, -3181, 1373, 9801),
                (0, 0, 0, 0, 0, 0, 0, 12207, -40371, -6040, 35631, 4626, 21024, -9218, -49),
                (0, 0, 0, 0, 0, 0, 0, 738, -7238, -8660, -119, 492, -3186, -837, 2313),
                (0, 0, 0, 0, 0, -41143, 0, 249, -26463, -4845, 26287, 8474, 30, -41143, -41143),
                (0, 0, 0, 0, 0, 0, 0, 1882, -63, 3828, -2899, -30126, 9190, 40811, 0),
                (0, 0, 0, 0, 0, 0, 0, 9059, -2220, 8099, -1236, 264, 3180, -7677, -876),
                (0, 0, 0, 0, 0, 0, 0, 20012, 127905, -7012, 2548, 56, -7776, -15932, 3213),
                (0, 0, 0, 0, 0, 0, 0, 15011, -7168, -285, -9449, 1145, -3299, 5914, -1165),
                (0, 0, 0, 0, 0, 0, 0, 4031, 241, 4351, -1454, -1849, 1438, 1637, -2727),
                (0, 0, 0, 0, 0, 0, 0, -110, 13472, -9559, -1012, 4271, -1974, 1907, -5062),
                (0, 0, 0, 0, 0, 0, 0, 48755, -23343, -6471, -142, -8312, 461, 4205, 240),
                (0, 0, 0, 0, 0, 0, 0, -3133, -12874, -10276, 1896, -120, -7060, -584, 2238),
                (0, 0, 0, 0, 0, 0, 0, -3066, 4400, -18769, 3062, -3023, 35020, -58653, 173),
                (0, 0, 0, 0, 0, 0, 0, 37, 7066, 1957, -8757, 3262, -5056, -10739, 15884),
                (0, 0, 0, 0, 0, 0, 0, -433, 722, 9770, 78, 402, -3111, -10631, 8010),
                (0, 0, 0, 0, 0, 0, 0, 5739, -120, 11913, 613, 9020, -7326, -6115, -792),
                (0, 0, 0, 0, 0, 0, 0, -5921, -231, 904, -13547, 3251, -1726, 846, -1895),
                (0, 0, 0, 0, 0, 0, 0, -3840, 2164, 1734, 17625, -10554, 5483, -808, 446),
                (0, 0, 0, 0, 0, 0, 0, -26930, 0, 19780, -8996, -1361, 14298, -9, -6768),
                (0, 0, 0, 0, 0, 0, 0, -87, 11574, -11205, -1285, 5541, -3762, -6195, 276),
                (0, 0, 0, 0, 0, 0, 0, 2043, -5541, 19454, -61046, -45828, 2170, -341, 512)
                );
    constant parent : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 4, 4, 5, 5, 6, 6, 3, 3),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 4, 4, 5, 5, 6, 6, 3, 3),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 6, 6, 5, 5),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 5, 5, 6, 6, 4, 4),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 6, 6, 5, 5),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6)
                );
    constant depth : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3)
                );
    constant iLeaf : intArray2D(nTrees-1 downto 0)(nLeaves-1 downto 0) := ((7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14)
                );
    constant value : tyArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := to_tyArray2D(value_int);
      constant threshold : txArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := to_txArray2D(threshold_int);
end Arrays0;