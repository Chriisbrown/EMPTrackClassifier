library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_misc.all;
  use ieee.numeric_std.all;

  use work.Constants.all;
  use work.Types.all;
  package Arrays0 is

    constant initPredict : ty := to_ty(0);
    constant feature : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((4, 1, 0, 0, 1, 2, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 4, 4, 4, 19, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 4, 4, 3, 17, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 1, 0, 3, 19, 2, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 1, 0, 0, 3, 2, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 4, 4, 4, 1, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 1, 0, 16, 17, 2, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 4, 4, 4, 1, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 4, 4, 3, 3, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 1, 0, 3, 3, 3, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 3, 2, 16, 17, 3, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 1, 4, 4, 0, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 1, 18, 3, 0, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 17, 2, 0, 3, 3, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 16, 0, 1, 3, 3, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 1, 4, 4, 0, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 19, 0, 1, 15, 3, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 1, 1, 4, 4, 3, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 4, 4, 10, -2, 17, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 1, 4, 3, 3, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 4, 4, 1, -2, 17, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 3, 18, 0, 1, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 4, 1, 0, -2, 0, 12, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 17, 2, 5, 3, 3, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 3, 2, 17, 16, 3, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 4, 1, 1, -2, 18, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 1, 4, 18, 4, 20, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 4, 0, 3, 17, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 4, 18, 0, -2, 18, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 18, 4, 18, 4, 16, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 16, 18, 17, 1, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 4, 0, 5, 16, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 18, 4, 18, 4, 16, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 16, 2, 20, 18, 16, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 16, 18, 17, 1, 7, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 17, 20, 7, 12, 12, 7, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 2, 18, 3, 5, 4, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 16, 2, 4, 20, 16, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 4, 1, 10, 0, 16, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 16, 18, 18, 1, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 18, 4, 4, 0, 17, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 16, 2, 20, 20, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (7, 17, 6, 5, 12, 20, 13, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 16, 2, 7, 18, 16, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 18, 4, 4, 3, 19, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 7, 18, 17, 13, 18, 20, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 7, 5, 17, 6, 8, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 1, 1, 2, -2, 5, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 17, 2, 7, 12, 20, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 18, 4, 4, 0, 17, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 7, 12, 17, 6, 5, 13, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 1, 18, 18, -2, 17, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 5, 17, 8, 0, 7, 13, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 18, 1, 18, -2, 5, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 17, 16, 7, 14, 17, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 17, 16, 7, 13, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 17, 8, 7, 12, 12, 9, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 18, 20, 4, 0, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 16, 17, 17, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 6, 17, 17, 7, 7, 12, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 16, 17, 16, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 3, 16, 5, -2, 4, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 18, 20, 18, 5, 19, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 18, 20, 4, 3, 17, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 18, 4, 18, 20, 18, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 5, 16, 8, 7, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 1, 16, 17, 17, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 17, 8, 7, 12, 17, 5, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 16, 6, 18, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 4, 18, 0, -2, 16, 20, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 7, 12, 5, 13, 5, 15, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 6, 16, 17, 7, 4, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 17, 8, 7, 12, 16, 9, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 5, 17, 18, 0, 6, 19, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 17, 2, 6, 14, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 20, 4, 10, 17, 18, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 2, 1, 17, -2, 3, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 6, 1, -2, -2, 17, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 18, 4, 4, 18, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 20, 18, 17, 2, 4, 20, -2, -2, -2, -2, -2, -2, -2, -2),
                (19, 6, 17, 17, 7, 20, 12, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 17, 16, 6, 14, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 3, 16, 17, 4, 8, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 19, -2, 7, 17, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 6, 17, -2, 5, 4, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 1, 4, 5, 17, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 18, 20, 4, 0, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (5, 8, 17, 17, 9, 4, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (19, 11, 12, 6, 16, 15, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 18, -2, 4, 3, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 17, 16, 7, 14, 4, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 3, 4, 18, 16, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 3, 5, -2, -2, 9, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 17, 16, 6, 17, 1, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 4, 18, 0, 0, 4, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 0, 4, 3, 16, 0, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 1, 4, 7, 16, 18, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (5, 8, 7, 17, 7, 12, 6, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 14, 0, 16, -2, 17, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 7, 14, 5, 13, 15, 13, -2, -2, -2, -2, -2, -2, -2, -2)
                );
    constant threshold_int : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((576, 258, 3012, 2482, 362, 2046, 3286, 0, 0, 0, 0, 0, 0, 0, 0),
                (304, 2780, 576, 576, 704, 320, 2094, 0, 0, 0, 0, 0, 0, 0, 0),
                (292, 2044, 576, 576, 1078, 412, 2616, 0, 0, 0, 0, 0, 0, 0, 0),
                (576, 204, 2924, 616, 320, 2046, 1242, 0, 0, 0, 0, 0, 0, 0, 0),
                (576, 226, 2892, 2348, 418, 2046, 1218, 0, 0, 0, 0, 0, 0, 0, 0),
                (318, 2046, 704, 576, 576, 502, 2656, 0, 0, 0, 0, 0, 0, 0, 0),
                (576, 180, 2846, 150, 412, 2046, 1290, 0, 0, 0, 0, 0, 0, 0, 0),
                (330, 2034, 704, 576, 576, 532, 2578, 0, 0, 0, 0, 0, 0, 0, 0),
                (280, 2034, 704, 576, 1058, 530, 2831, 0, 0, 0, 0, 0, 0, 0, 0),
                (576, 170, 2066, 512, 420, 1328, 1194, 0, 0, 0, 0, 0, 0, 0, 0),
                (576, 540, 2046, 198, 514, 1382, 3018, 0, 0, 0, 0, 0, 0, 0, 0),
                (264, 1956, 522, 576, 704, 1816, 310, 0, 0, 0, 0, 0, 0, 0, 0),
                (240, 1820, 474, 1361, 1184, 2208, 302, 0, 0, 0, 0, 0, 0, 0, 0),
                (576, 394, 2046, 926, 718, 1382, 2930, 0, 0, 0, 0, 0, 0, 0, 0),
                (576, 220, 2074, 130, 630, 1312, 208, 0, 0, 0, 0, 0, 0, 0, 0),
                (362, 1638, 640, 576, 704, 2312, 336, 0, 0, 0, 0, 0, 0, 0, 0),
                (576, 320, 2068, 132, 64, 1311, 2754, 0, 0, 0, 0, 0, 0, 0, 0),
                (1544, 394, 212, 576, 576, 1390, 264, 0, 0, 0, 0, 0, 0, 0, 0),
                (1438, 576, 704, 64, 0, 412, 1512, 0, 0, 0, 0, 0, 0, -256, -256),
                (390, 1368, 644, 576, 866, 646, 344, 0, 0, 0, 0, 0, 0, 0, 0),
                (1386, 576, 704, 250, 0, 392, 1410, 0, 0, 0, 0, 0, 0, -256, -256),
                (198, 1546, 680, 1294, 2748, 574, 704, 0, 0, 0, 0, 0, 0, 0, 0),
                (1278, 576, 152, 512, 0, 2566, 64, 0, 0, 0, 0, 0, 0, -256, -256),
                (576, 116, 2046, 64, 438, 1388, 152, 0, 0, 0, 0, 0, 0, 0, 0),
                (704, 660, 2044, 450, 192, 1382, 3578, 0, 0, 0, 0, 0, 0, 0, 0),
                (1298, 576, 446, 146, 0, -1128, 666, 0, 0, 0, 0, 0, 0, -256, -256),
                (1040, 386, 704, 1248, 576, 192, 1657, 0, 0, 0, 0, 0, 0, 0, 0),
                (140, 2188, 704, 742, 1228, 124, 2022, 0, 0, 0, 0, 0, 0, 0, 0),
                (1138, 576, 1084, 456, 0, -964, 704, 0, 0, 0, 0, 0, 0, -256, -256),
                (874, 1234, 704, -1151, 704, 242, 3578, 0, 0, 0, 0, 0, 0, 0, 0),
                (570, 926, 302, 1196, 404, 762, 0, 0, 0, 0, 0, 0, 0, -256, -256),
                (138, 2188, 704, 730, 64, 176, 2626, 0, 0, 0, 0, 0, 0, 0, 0),
                (866, 1241, 576, -1271, 576, 268, 1574, 0, 0, 0, 0, 0, 0, 0, 0),
                (704, 130, 2044, 576, 986, 184, 3699, 0, 0, 0, 0, 0, 0, 0, 0),
                (532, 920, 292, -1061, 396, 770, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (860, 456, 576, 64, 64, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (124, 2042, -1038, 1036, 64, 704, 1218, 0, 0, 0, 0, 0, 0, 0, 0),
                (704, 138, 2044, 576, 192, 200, 3696, 0, 0, 0, 0, 0, 0, 0, 0),
                (2448, 576, 106, 64, 866, 68, 704, 0, 0, 0, 0, 0, 0, 0, 0),
                (570, 712, 300, 1211, -1338, 764, 0, 0, 0, 0, 0, 0, 0, -256, -256),
                (1241, -971, 704, 576, 2448, 602, 0, 0, 0, 0, 0, 0, 0, -256, -256),
                (602, 774, 284, 240, 192, 704, 430, 0, 0, 0, 0, 0, 0, 0, 0),
                (64, 294, 64, 64, 64, 576, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (704, 138, 2042, 64, -1114, 186, 3076, 0, 0, 0, 0, 0, 0, 0, 0),
                (806, -731, 576, 576, 712, 320, 2017, 0, 0, 0, 0, 0, 0, 0, 0),
                (122, 64, 784, 284, 64, -1346, 576, 0, 0, 0, 0, 0, 0, 0, 0),
                (2284, 64, 64, 284, 64, 64, 704, 0, 0, 0, 0, 0, 0, 0, 0),
                (686, 360, 644, 192, 0, 64, 344, 0, 0, 0, 0, 0, 0, -256, -256),
                (948, 534, 972, 64, 64, 704, 192, 0, 0, 0, 0, 0, 0, 0, 0),
                (1414, -941, 704, 576, 2486, 602, 0, 0, 0, 0, 0, 0, 0, -256, -256),
                (390, 64, 64, 296, 64, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (496, 582, 941, 1084, 0, 390, 704, 0, 0, 0, 0, 0, 0, -256, -256),
                (98, 64, 392, 64, 1650, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (550, 881, 756, -941, 0, 64, 356, 0, 0, 0, 0, 0, 0, -256, -256),
                (2036, 556, 344, 64, 64, 678, 0, 0, 0, 0, 0, 0, 0, -256, -256),
                (1560, 384, 360, 64, 64, 0, 0, 0, 0, 0, 0, -256, -256, -256, -256),
                (656, 284, 64, 64, 64, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (1421, -836, 576, 576, 2284, 0, 0, 0, 0, 0, 0, -256, -256, -256, -256),
                (764, 574, 302, 92, 282, 0, 0, 0, 0, 0, 0, -256, -256, -256, -256),
                (686, 64, 268, 134, 64, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (814, 774, 366, 74, 112, 0, 0, 0, 0, 0, 0, -256, -256, -256, -256),
                (104, 1292, 180, 64, 0, 704, 92, 0, 0, 0, 0, 0, 0, -256, -256),
                (656, -731, 576, -1541, 64, 320, 0, 0, 0, 0, 0, 0, 0, -256, -256),
                (1398, -1346, 576, 576, 2042, 604, 0, 0, 0, 0, 0, 0, 0, -256, -256),
                (370, 828, 576, -566, 576, 994, 0, 0, 0, 0, 0, 0, 0, -256, -256),
                (850, 64, 364, 64, 64, 0, 0, 0, 0, 0, 0, -256, -256, -256, -256),
                (886, 68, 342, 186, 282, 0, 0, 0, 0, 0, 0, -256, -256, -256, -256),
                (660, 282, 64, 64, 64, 280, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (908, 516, 366, 64, 1548, 0, 0, 0, 0, 0, 0, -256, -256, -256, -256),
                (-1338, 576, 626, 3861, 0, 108, 576, 0, 0, 0, 0, 0, 0, -256, -256),
                (296, 64, 64, 64, 64, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (2176, 64, 112, 122, 64, 704, 268, 0, 0, 0, 0, 0, 0, 0, 0),
                (660, 294, 64, 64, 64, 168, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (72, 64, 104, -1001, 2154, 64, 192, 0, 0, 0, 0, 0, 0, 0, 0),
                (954, 552, 838, 64, 64, 364, 100, 0, 0, 0, 0, 0, 0, 0, 0),
                (360, 576, 576, 64, 186, -1144, 0, 0, 0, 0, 0, 0, 0, -256, -256),
                (564, 192, 102, 42, 0, 1390, 300, 0, 0, 0, 0, 0, 0, -256, -256),
                (492, 64, 956, 0, 0, 556, 0, 0, 0, -256, -256, -256, -256, -256, -256),
                (368, -1338, 576, 704, 626, 0, 0, 0, 0, 0, 0, -256, -256, -256, -256),
                (-566, 576, 626, 304, 1976, 576, 576, 0, 0, 0, 0, 0, 0, 0, 0),
                (192, 64, 262, 136, 64, 320, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (2042, 554, 240, 64, 64, 0, 0, 0, 0, 0, 0, -256, -256, -256, -256),
                (2286, 878, 98, 62, 704, 64, 576, 0, 0, 0, 0, 0, 0, 0, 0),
                (916, 192, 0, 64, 246, 0, 0, 0, 0, -256, -256, -256, -256, -256, -256),
                (70, 64, 78, 0, 64, 704, 184, 0, 0, 0, 0, 0, 0, -256, -256),
                (370, 68, 576, 64, 92, 0, 0, 0, 0, 0, 0, -256, -256, -256, -256),
                (1458, -1451, 576, 576, 732, 0, 0, 0, 0, 0, 0, -256, -256, -256, -256),
                (64, 64, 92, 246, 64, 704, 576, 0, 0, 0, 0, 0, 0, 0, 0),
                (192, 64, 64, 64, 98, 64, 266, 0, 0, 0, 0, 0, 0, 0, 0),
                (1548, -566, 0, 704, 986, 0, 0, 0, 0, -256, -256, -256, -256, -256, -256),
                (2450, 312, 110, 64, 64, 704, 96, 0, 0, 0, 0, 0, 0, 0, 0),
                (370, 2042, 576, -1541, 240, 0, 0, 0, 0, 0, 0, -256, -256, -256, -256),
                (70, 1048, 64, 0, 0, 64, 116, 0, 0, 0, 0, -256, -256, -256, -256),
                (68, 180, 360, 64, 244, 822, 576, 0, 0, 0, 0, 0, 0, 0, 0),
                (-686, 704, 618, 3600, 2596, 576, 576, 0, 0, 0, 0, 0, 0, 0, 0),
                (1391, 2448, 576, 1304, 68, 2844, 0, 0, 0, 0, 0, 0, 0, -256, -256),
                (360, 850, 576, 64, 316, 814, 1394, 0, 0, 0, 0, 0, 0, 0, 0),
                (64, 64, 64, 262, 64, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0),
                (68, 64, 2344, 296, 0, 72, 68, 0, 0, 0, 0, 0, 0, -256, -256),
                (282, 64, 64, 64, 64, 64, 64, 0, 0, 0, 0, 0, 0, 0, 0)
                );
    constant children_left : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 13, 9, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 13, 9, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 13, 9, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 13, 9, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 13, 9, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 13, 9, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 13, 9, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 13, 9, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 13, 9, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 13, 9, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 13, 9, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 9, 11, 7, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 9, 5, 7, -1, -1, -1, -1, 11, 13, -1, -1, -1, -1),
                (1, 3, 5, 13, 7, 9, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 9, 5, 7, -1, -1, -1, -1, 11, 13, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 11, 13, 7, 9, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 13, 9, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1)
                );
    constant children_right : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 14, 10, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 14, 10, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 14, 10, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 14, 10, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 14, 10, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 14, 10, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 14, 10, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 14, 10, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 14, 10, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 14, 10, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 14, 10, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 10, 12, 8, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 10, 6, 8, -1, -1, -1, -1, 12, 14, -1, -1, -1, -1),
                (2, 4, 6, 14, 8, 10, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 10, 6, 8, -1, -1, -1, -1, 12, 14, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 12, 14, 8, 10, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 14, 10, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1)
                );
    constant value_int : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((0, 0, 0, 0, 0, 0, 0, 14, -10, -12, -24, 27, 19, 3, -13),
                (0, 0, 0, 0, 0, 0, 0, 9, 23, -10, 8, -22, -9, 22, -5),
                (0, 0, 0, 0, 0, 0, 0, 16, 23, 12, -10, -20, -7, 14, -11),
                (0, 0, 0, 0, 0, 0, 0, 12, -8, -17, -1, 21, 14, 4, -10),
                (0, 0, 0, 0, 0, 0, 0, 11, -5, -8, -18, 20, 13, 5, -8),
                (0, 0, 0, 0, 0, 0, 0, 13, 19, -2, 11, -8, -18, 15, 0),
                (0, 0, 0, 0, 0, 0, 0, -5, 11, -14, 1, 18, 11, 3, -9),
                (0, 0, 0, 0, 0, 0, 0, 12, 17, -2, 10, -7, -16, 13, 0),
                (0, 0, 0, 0, 0, 0, 0, 11, 17, 8, -8, -5, -15, 13, -1),
                (0, 0, 0, 0, 0, 0, 0, 10, -4, -3, -14, 16, 0, 9, -7),
                (0, 0, 0, 0, 0, 0, 0, -7, 8, -13, 0, 16, -3, 8, -5),
                (0, 0, 0, 0, 0, 0, 0, 10, 15, 1, 10, 9, -6, -15, -3),
                (0, 0, 0, 0, 0, 0, 0, 14, 0, 6, -7, 6, -6, -13, -3),
                (0, 0, 0, 0, 0, 0, 0, 8, -9, 13, -5, 14, -3, 7, -4),
                (0, 0, 0, 0, 0, 0, 0, 0, -11, 6, -6, 14, 0, 7, -2),
                (0, 0, 0, 0, 0, 0, 0, 8, 14, 0, 8, 0, -9, -14, 0),
                (0, 0, 0, 0, 0, 0, 0, 2, -8, 13, -1, 13, 0, 6, -3),
                (0, 0, 0, 0, 0, 0, 0, 8, 13, -7, 10, 5, -7, -9, 0),
                (0, 0, 0, 0, 13, 0, 0, 7, -9, -5, 6, 8, -6, 13, 13),
                (0, 0, 0, 0, 0, 0, 0, 7, 13, 4, -4, -1, -9, -13, 0),
                (0, 0, 0, 0, 12, 0, 0, 8, -3, -5, 5, 8, -4, 12, 12),
                (0, 0, 0, 0, 0, 0, 0, 11, 0, 5, -2, 2, -9, -10, 1),
                (0, 0, 0, 0, 12, 0, 0, 10, 0, 6, 0, -7, 1, 12, 12),
                (0, 0, 0, 0, 0, 0, 0, 0, -12, 5, -4, 11, -1, 4, -1),
                (0, 0, 0, 0, 0, 0, 0, 0, 11, -10, -3, 11, 0, 5, -5),
                (0, 0, 0, 0, 11, 0, 0, 9, 0, -11, 2, -5, -12, 11, 11),
                (0, 0, 0, 0, 0, 0, 0, 10, 0, -3, 7, 6, -4, 6, -6),
                (0, 0, 0, 0, 0, 0, 0, 11, 7, 3, -3, -9, -1, 10, 2),
                (0, 0, 0, 0, 11, 0, 0, 9, 0, -9, 2, -13, 1, 11, 11),
                (0, 0, 0, 0, 0, 0, 0, -10, 4, -14, 1, -9, -2, 2, -4),
                (0, 0, 0, 0, 0, 0, 0, 9, 0, -1, 5, -7, -13, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, 10, 6, 6, 1, -7, 0, 7, -1),
                (0, 0, 0, 0, 0, 0, 0, -11, 3, -14, 0, -9, -1, 0, -4),
                (0, 0, 0, 0, 0, 0, 0, -8, 0, 2, -9, 12, 6, 3, -5),
                (0, 0, 0, 0, 0, 0, 0, 0, 8, -1, 5, -6, -12, -3, 1),
                (0, 0, 0, 0, 0, 0, 0, -6, 4, -5, 9, -9, -3, -9, 1),
                (0, 0, 0, 0, 0, 0, 0, 7, 0, 6, 0, -10, 0, 0, -11),
                (0, 0, 0, 0, 0, 0, 0, -8, -1, 6, -1, 11, 5, 2, -5),
                (0, 0, 0, 0, 0, 0, 0, 1, -12, 9, 3, -2, 2, -5, 0),
                (0, 0, 0, 0, 0, 0, 0, 8, 0, -10, 1, -5, -11, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, -10, 0, 3, -1, -11, 0, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, 8, 2, 4, -1, -9, 0, 0, -4),
                (0, 0, 0, 0, 0, 0, 0, 4, -18, -10, 4, -10, 0, 5, -3),
                (0, 0, 0, 0, 0, 0, 0, -8, -2, -8, 1, 11, 3, 2, -2),
                (0, 0, 0, 0, 0, 0, 0, -6, 0, 3, -1, -9, 0, 3, -2),
                (0, 0, 0, 0, 0, 0, 0, -14, 3, 5, -1, -9, 0, -7, 0),
                (0, 0, 0, 0, 0, 0, 0, -14, 4, -8, 5, 0, 8, -4, 0),
                (0, 0, 0, 0, 0, 0, 0, 8, 2, 3, -1, -8, 0, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, -3, 3, -2, 8, -8, 0, -4, 0),
                (0, 0, 0, 0, 0, 0, 0, -7, 0, 2, -1, -11, 0, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, -13, 0, -7, 2, 0, -13, -8, 6),
                (0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 3, -6, 2, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, 2, 10, 4, 0, -7, 0, -8, 3),
                (0, 0, 0, 0, 0, 0, 0, 0, 7, 2, -1, -8, 0, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, -3, 1, 10, 3, -6, 0, 0, 0),
                (0, 0, 0, 0, 0, -5, 3, -5, 2, -8, 5, -5, -5, 3, 3),
                (0, 0, 0, 0, 0, 0, 0, -12, 2, -7, 5, -8, -2, -4, 1),
                (0, 0, 0, 0, 0, -9, 0, -5, 0, 2, 0, -9, -9, 0, 0),
                (0, 0, 0, 0, 0, -9, 0, 0, 7, -1, 1, -9, -9, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, -6, 2, 1, 7, -10, 0, -7, 2),
                (0, 0, 0, 0, 0, -8, 0, 0, 5, -2, 1, -8, -8, 0, 0),
                (0, 0, 0, 0, -1, 0, 0, 5, 2, -4, 2, -3, 1, -1, -1),
                (0, 0, 0, 0, 0, 0, 1, -8, -1, 4, 1, -5, 0, 1, 1),
                (0, 0, 0, 0, 0, 0, 0, -8, 0, 1, -3, -8, 0, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, -2, 1, -4, 0, 11, 0, 0, 0),
                (0, 0, 0, 0, 0, -8, 0, 0, 8, -2, 1, -8, -8, 0, 0),
                (0, 0, 0, 0, 0, -9, 0, 4, 1, -1, 1, -9, -9, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, -10, 1, -5, 4, -6, -2, 5, 0),
                (0, 0, 0, 0, 0, -8, 0, 0, 5, 0, -8, -8, -8, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, -7, 0, -1, 1, -3, 1, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, 12, -11, 1, -5, 5, -7, 5, -1),
                (0, 0, 0, 0, 0, 0, 0, -10, 1, -1, 4, -5, 1, -1, 1),
                (0, 0, 0, 0, 0, 0, 0, -7, 1, -4, 3, -5, -1, -2, 2),
                (0, 0, 0, 0, 0, 0, 0, 0, 5, 3, 0, -9, 0, 3, -1),
                (0, 0, 0, 0, 0, 0, 0, -5, 1, 9, 2, -6, 0, -4, 0),
                (0, 0, 0, 0, 0, 0, 0, 0, -8, 2, -6, 0, 7, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, 0, 6, 1, -1, -1, 0, 0, 0),
                (0, 0, 0, 0, 5, 0, -7, 0, 2, 0, 0, 5, 5, -7, -7),
                (0, 0, 0, 0, 0, 8, 0, -6, 0, 0, -2, 8, 8, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, -3, 0, 3, -1, 2, 0, -2, 1),
                (0, 0, 0, 0, 0, 0, 0, -7, 0, -5, 3, -8, -2, -5, 1),
                (0, 0, 0, 0, 0, -5, 0, -3, 0, 7, 1, -5, -5, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, -1, 1, -5, 0, -5, 0, 1, -1),
                (0, 0, -6, 0, 0, -5, 2, -5, 0, -6, -6, -6, -6, -6, -6),
                (0, 0, 0, 0, 0, 0, 0, 0, 8, -3, 2, 2, 0, 0, 0),
                (0, 0, 0, 0, 0, 7, 0, 3, 1, -2, 0, 7, 7, 0, 0),
                (0, 0, 0, 0, 0, -6, 0, -6, 0, 2, 0, -6, -6, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, -7, 1, -6, 8, -5, 2, 2, -1),
                (0, 0, 0, 0, 0, 0, 0, -4, 1, 0, 11, -9, 0, -3, 1),
                (0, 0, -6, 0, 0, -2, 0, 1, -1, -6, -6, -6, -6, -6, -6),
                (0, 0, 0, 0, 0, 0, 0, -5, 1, 6, 0, -5, 0, 1, -1),
                (0, 0, 0, 0, 0, 6, 0, -5, 0, -4, 0, 6, 6, 0, 0),
                (0, 0, 0, 5, 0, 0, 0, -1, 6, -2, 0, 5, 5, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, 0, 3, -1, 1, 0, -4, 6, -1),
                (0, 0, 0, 0, 0, 0, 0, -2, 0, 2, -1, 1, 0, -2, 0),
                (0, 0, 0, 0, 0, 0, 0, 1, -4, -3, 0, -7, 0, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, -1, 0, -6, 0, 6, 0, -2, 0),
                (0, 0, 0, 0, 0, 0, 0, -5, 1, 19, 3, -7, 1, -3, 1),
                (0, 0, 0, 0, 0, 0, 0, 2, 0, -1, 1, -3, 0, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, 13, -8, 1, -4, 5, -4, -7, 0)
                );
    constant parent : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 5, 5, 6, 6, 4, 4),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 5, 5, 6, 6, 4, 4),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 5, 5, 6, 6, 4, 4),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 5, 5, 6, 6, 4, 4),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 5, 5, 6, 6, 4, 4),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 5, 5, 6, 6, 4, 4),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 5, 5, 6, 6, 4, 4),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 5, 5, 6, 6, 4, 4),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 5, 5, 6, 6, 4, 4),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 5, 5, 6, 6, 4, 4),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 5, 5, 6, 6, 4, 4),
                (-1, 0, 0, 1, 1, 2, 2, 5, 5, 3, 3, 4, 4, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 3, 3, 4, 4, 2, 2, 9, 9, 10, 10),
                (-1, 0, 0, 1, 1, 2, 2, 4, 4, 5, 5, 6, 6, 3, 3),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 3, 3, 4, 4, 2, 2, 9, 9, 10, 10),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 5, 5, 6, 6, 3, 3, 4, 4),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 5, 5, 6, 6, 4, 4),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6)
                );
    constant depth : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 3, 3, 3, 3, 2, 2, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 3, 3, 3, 3, 2, 2, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3)
                );
    constant iLeaf : intArray2D(nTrees-1 downto 0)(nLeaves-1 downto 0) := ((7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (5, 6, 7, 8, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (5, 6, 7, 8, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14)
                );
    constant value : tyArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := to_tyArray2D(value_int);
      constant threshold : txArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := to_txArray2D(threshold_int);
end Arrays0;