library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_misc.all;
  use ieee.numeric_std.all;

  use work.Constants.all;
  use work.Types.all;
  package Arrays0 is

    constant initPredict : ty := to_ty(0);
    constant feature : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((4, 3, 0, 2, 3, 0, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 3, 0, 0, 3, 2, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 3, 0, 2, 19, 0, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 0, 4, 4, 4, 3, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 3, 0, 16, 19, 0, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 0, 4, 18, 2, 2, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 19, 0, 0, 2, 2, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 0, 3, 18, 4, 0, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 0, 3, 2, 0, 2, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 18, 0, 16, 17, 1, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 0, 3, 18, 17, 2, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 18, 4, 0, 4, 17, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 0, 17, 1, 4, 4, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 17, 4, 7, 15, 12, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 2, 4, 0, 16, 17, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 2, 4, 17, 4, 12, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 4, 3, 17, 16, 18, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 5, 17, 9, 4, 4, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 3, 16, 0, 16, 20, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 2, 4, 17, 16, 12, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 18, 3, 2, 4, 16, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 5, 17, 9, 20, 7, 12, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 2, 17, 7, 20, 7, 12, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 0, 16, 1, 5, 3, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 2, 4, 0, 16, 17, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (20, 17, 16, 5, 2, 0, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 5, 4, 9, 1, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 17, 16, 7, 14, 19, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 20, 16, 13, 6, 20, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 2, 4, 17, 12, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (20, 17, 16, 5, 2, 0, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 5, 1, 8, 16, 20, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (7, 12, 6, 5, 13, 4, 19, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 3, 0, 7, 16, 16, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 2, 18, 7, 20, 17, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 17, 20, 7, 19, 10, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 0, 16, 1, 0, 3, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 18, 16, 7, 4, 20, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 7, 12, 5, 19, 17, 15, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 6, 19, 4, 7, 7, 12, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 3, 4, 17, 16, 3, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 17, 8, 6, 19, 20, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 16, 4, 1, 2, 3, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 20, 16, 17, 1, 1, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 18, 17, 2, 3, 3, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 17, 16, 7, 14, 19, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 17, 16, 6, 2, 4, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 16, 2, 3, 0, 0, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 16, 2, 0, 4, 17, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 2, 4, 18, 4, 18, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 0, 19, 16, 16, 6, 12, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 7, 14, 5, 13, 15, 13, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 4, 5, 16, 16, 9, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (11, 8, 15, 5, 7, 17, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (11, 1, 15, 16, 19, 4, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 0, 3, 4, 5, 5, 14, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 18, 10, 17, 3, 11, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 0, 2, 4, 1, 1, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 5, 16, 17, 9, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 4, 2, 16, 16, 17, 8, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 20, 14, 8, 6, 16, 19, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 17, 3, 20, 14, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 0, 17, 16, 0, 7, 14, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 17, 11, 18, 16, 8, 19, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 2, 16, 17, 8, -2, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 3, 0, 16, 3, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 1, 16, 12, 1, 14, 15, -2, -2, -2, -2, -2, -2, -2, -2),
                (5, 16, 16, 1, 9, 4, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 7, 13, 4, 6, 17, 12, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 16, 10, 17, 4, 4, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 16, 4, 3, 16, 3, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 16, 16, 4, 4, 17, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 3, 18, 3, 16, 3, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 1, 19, 16, 16, 16, 12, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 16, 2, 0, 1, 2, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 8, 16, 10, 5, 20, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 18, 16, 16, 20, 19, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 13, 13, 17, 4, 17, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 3, 17, 16, 16, 0, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 3, 16, 9, 16, 0, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 4, 18, 0, 2, 5, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 13, 13, 17, 19, 20, 15, -2, -2, -2, -2, -2, -2, -2, -2),
                (8, 10, 20, 19, 0, 3, 6, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 16, 16, 4, 4, 4, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, -2, 3, 16, 3, -2, -2, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 3, 2, 5, 16, 0, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 1, 4, 16, 16, 19, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 4, 0, 16, 16, 17, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (20, 17, 17, 6, 7, 6, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 3, 2, 16, 16, 18, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 20, 16, 2, 17, 0, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 5, 1, 16, 16, 5, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 0, 2, 18, 0, 3, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 5, 16, 9, 9, 19, 20, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 4, 19, 10, 16, 17, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 16, 17, 0, 8, 20, 12, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 5, 5, 14, 16, 9, 9, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 1, 16, 0, 16, -2, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 1, 19, 4, 16, 17, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 2, 14, 3, 17, 4, 0, -2, -2, -2, -2, -2, -2, -2, -2)
                );
    constant threshold_int : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((288, 30, 215, 92, 64, 174, 129, 0, 0, 0, 0, 0, 0, 0, 0),
                (288, 24, 227, 171, 58, 148, 122, 0, 0, 0, 0, 0, 0, 0, 0),
                (288, 42, 202, 79, 160, 154, 138, 0, 0, 0, 0, 0, 0, 0, 0),
                (44, 196, 352, 288, 352, 71, 265, 0, 0, 0, 0, 0, 0, 0, 0),
                (288, 11, 261, 89, 160, 167, 34, 0, 0, 0, 0, 0, 0, 0, 0),
                (52, 181, 352, 707, 116, 81, 194, 0, 0, 0, 0, 0, 0, 0, 0),
                (288, 160, 292, 112, 102, 135, 99, 0, 0, 0, 0, 0, 0, 0, 0),
                (58, 153, 90, 632, 352, 146, 160, 0, 0, 0, 0, 0, 0, 0, 0),
                (35, 272, 80, 135, 358, 102, 108, 0, 0, 0, 0, 0, 0, 0, 0),
                (288, 467, 159, 97, 263, 77, 153, 0, 0, 0, 0, 0, 0, 0, 0),
                (69, 145, 99, 729, 198, 98, 154, 0, 0, 0, 0, 0, 0, 0, 0),
                (113, 572, 352, 315, 352, 259, 159, 0, 0, 0, 0, 0, 0, 0, 0),
                (72, 130, 64, 27, 352, 352, 50, 0, 0, 0, 0, 0, 0, 0, 0),
                (125, 222, 288, 32, 32, 32, 309, 0, 0, 0, 0, 0, 0, 0, 0),
                (9, 148, 352, 369, 122, 63, 199, 0, 0, 0, 0, 0, 0, 0, 0),
                (542, 101, 288, 197, 352, 32, 139, 0, 0, 0, 0, 0, 0, 0, 0),
                (133, 288, 90, 59, 117, 669, 111, 0, 0, 0, 0, 0, 0, 0, 0),
                (2, 32, 277, 32, 352, 352, 146, 0, 0, 0, 0, 0, 0, 0, 0),
                (327, 100, 14, 109, 154, 352, 379, 0, 0, 0, 0, 0, 0, 0, 0),
                (426, 154, 288, 271, 111, 32, 149, 0, 0, 0, 0, 0, 0, 0, 0),
                (364, 688, 0, 98, 352, 10, 77, 0, 0, 0, 0, 0, 0, 0, 0),
                (-17, 32, 194, 32, 352, 32, 32, 0, 0, 0, 0, 0, 0, 0, 0),
                (49, 140, 136, 32, 288, 32, 32, 0, 0, 0, 0, 0, 0, 0, 0),
                (109, 104, 128, -11, 32, 124, 136, 0, 0, 0, 0, 0, 0, 0, 0),
                (729, 153, 352, 368, 125, 263, 182, 0, 0, 0, 0, 0, 0, 0, 0),
                (352, 51, 69, 32, 74, 339, 68, 0, 0, 0, 0, 0, 0, 0, 0),
                (347, 32, 288, 32, 60, 79, 127, 0, 0, 0, 0, 0, 0, 0, 0),
                (121, 262, 139, 32, 32, 224, 135, 0, 0, 0, 0, 0, 0, 0, 0),
                (302, 96, 10, 32, 32, 352, 68, 0, 0, 0, 0, 0, 0, 0, 0),
                (362, 165, 288, 137, 32, 120, 22, 0, 0, 0, 0, 0, 0, 0, 0),
                (352, 47, 96, 32, 64, 320, 236, 0, 0, 0, 0, 0, 0, 0, 0),
                (-42, 32, 27, 32, 114, 288, 139, 0, 0, 0, 0, 0, 0, 0, 0),
                (32, 32, 32, 32, 32, 288, 96, 0, 0, 0, 0, 0, 0, 0, 0),
                (391, 113, 419, 32, 118, 12, 90, 0, 0, 0, 0, 0, 0, 0, 0),
                (-20, 140, 771, 32, 288, 136, 887, 0, 0, 0, 0, 0, 0, 0, 0),
                (21, 60, 288, 32, 96, 32, 83, 0, 0, 0, 0, 0, 0, 0, 0),
                (121, 80, 123, -67, 398, 126, 15, 0, 0, 0, 0, 0, 0, 0, 0),
                (182, 816, 179, 32, 352, 288, 306, 0, 0, 0, 0, 0, 0, 0, 0),
                (146, 32, 32, 32, 96, 161, 32, 0, 0, 0, 0, 0, 0, 0, 0),
                (46, 32, 96, 288, 32, 32, 32, 0, 0, 0, 0, 0, 0, 0, 0),
                (187, 129, 288, 152, 139, 60, 12, 0, 0, 0, 0, 0, 0, 0, 0),
                (110, 68, 32, 32, 96, 96, 216, 0, 0, 0, 0, 0, 0, 0, 0),
                (186, 2, 288, 185, 180, 56, -64, 0, 0, 0, 0, 0, 0, 0, 0),
                (-4, 288, 2, 24, -67, 164, 137, 0, 0, 0, 0, 0, 0, 0, 0),
                (416, 309, 90, -28, -87, -57, 67, 0, 0, 0, 0, 0, 0, 0, 0),
                (130, 279, 122, 32, 32, 224, 6, 0, 0, 0, 0, 0, 0, 0, 0),
                (-35, 93, 154, 32, 21, 288, 288, 0, 0, 0, 0, 0, 0, 0, 0),
                (819, 1, 221, 24, 379, 173, 0, 0, 0, 0, 0, 0, 0, -128, -128),
                (-37, 107, 63, 204, 352, 133, 352, 0, 0, 0, 0, 0, 0, 0, 0),
                (186, 224, 288, 857, 352, 572, 90, 0, 0, 0, 0, 0, 0, 0, 0),
                (67, 212, 96, 21, 111, 32, 32, 0, 0, 0, 0, 0, 0, 0, 0),
                (151, 32, 32, 32, 32, 32, 32, 0, 0, 0, 0, 0, 0, 0, 0),
                (68, 288, 32, 185, 38, 32, 124, 0, 0, 0, 0, 0, 0, 0, 0),
                (32, 32, 32, 32, 32, 126, 288, 0, 0, 0, 0, 0, 0, 0, 0),
                (32, 235, 32, 14, 160, 288, 288, 0, 0, 0, 0, 0, 0, 0, 0),
                (3, 203, 138, 288, 32, 32, 32, 0, 0, 0, 0, 0, 0, 0, 0),
                (420, 302, 32, 68, 91, 32, -21, 0, 0, 0, 0, 0, 0, 0, 0),
                (3, 197, 224, 288, 219, 433, 143, 0, 0, 0, 0, 0, 0, 0, 0),
                (27, 132, 32, 17, 157, 32, 142, 0, 0, 0, 0, 0, 0, 0, 0),
                (15, 288, 80, 38, 94, 124, 32, 0, 0, 0, 0, 0, 0, 0, 0),
                (134, 160, 32, 32, 32, 72, 160, 0, 0, 0, 0, 0, 0, 0, 0),
                (-34, 125, -12, 160, 32, 92, 186, 0, 0, 0, 0, 0, 0, 0, 0),
                (3, 203, 161, 2, 264, 32, 32, 0, 0, 0, 0, 0, 0, 0, 0),
                (44, 17, 32, 144, 107, 32, 96, 0, 0, 0, 0, 0, 0, 0, 0),
                (143, 106, 104, 122, 32, 0, 155, 0, 0, 0, 0, 0, 0, -128, -128),
                (-204, 53, 391, 72, 84, 8, 14, 0, 0, 0, 0, 0, 0, 0, 0),
                (124, -64, 140, 32, -63, 32, 32, 0, 0, 0, 0, 0, 0, 0, 0),
                (32, 65, 130, 244, 32, 352, 288, 0, 0, 0, 0, 0, 0, 0, 0),
                (158, 32, 32, 288, 32, 185, 32, 0, 0, 0, 0, 0, 0, 0, 0),
                (71, 16, 32, 45, 288, 288, 288, 0, 0, 0, 0, 0, 0, 0, 0),
                (187, 2, 352, 21, 165, 80, 187, 0, 0, 0, 0, 0, 0, 0, 0),
                (330, 16, 32, 288, 288, 211, 154, 0, 0, 0, 0, 0, 0, 0, 0),
                (-67, -68, 857, -69, 162, 44, 217, 0, 0, 0, 0, 0, 0, 0, 0),
                (66, 232, 96, 14, 125, 58, 32, 0, 0, 0, 0, 0, 0, 0, 0),
                (432, 3, 102, 200, -47, 98, 119, 0, 0, 0, 0, 0, 0, 0, 0),
                (127, 32, 171, 32, 32, 32, 139, 0, 0, 0, 0, 0, 0, 0, 0),
                (182, 763, 111, 3, 96, 288, 352, 0, 0, 0, 0, 0, 0, 0, 0),
                (157, 32, 32, 128, 352, 184, 196, 0, 0, 0, 0, 0, 0, 0, 0),
                (187, 141, 161, 165, 104, 169, 206, 0, 0, 0, 0, 0, 0, 0, 0),
                (-42, 52, 9, 32, 83, 225, 192, 0, 0, 0, 0, 0, 0, 0, 0),
                (51, 288, 317, 73, 66, 32, 97, 0, 0, 0, 0, 0, 0, 0, 0),
                (186, 32, 32, 129, 160, 32, 32, 0, 0, 0, 0, 0, 0, 0, 0),
                (32, 32, 160, 96, 209, 23, 32, 0, 0, 0, 0, 0, 0, 0, 0),
                (52, 142, 91, 288, 288, 352, 168, 0, 0, 0, 0, 0, 0, 0, 0),
                (1, 0, -17, 92, 35, 0, 0, 0, 0, -128, -128, -128, -128, -128, -128),
                (416, 104, 14, 32, 138, 425, 34, 0, 0, 0, 0, 0, 0, 0, 0),
                (186, 189, 288, 29, 49, 160, 76, 0, 0, 0, 0, 0, 0, 0, 0),
                (79, 288, 142, 143, 36, 92, 46, 0, 0, 0, 0, 0, 0, 0, 0),
                (160, 135, 145, 32, 32, 32, 245, 0, 0, 0, 0, 0, 0, 0, 0),
                (115, 51, 5, 108, 122, 399, 174, 0, 0, 0, 0, 0, 0, 0, 0),
                (-45, 288, 186, -8, 66, 416, 352, 0, 0, 0, 0, 0, 0, 0, 0),
                (267, 32, 220, 88, 111, 32, 212, 0, 0, 0, 0, 0, 0, 0, 0),
                (-87, 350, -158, 444, 359, 57, 272, 0, 0, 0, 0, 0, 0, 0, 0),
                (179, 32, 113, 32, 32, 288, 288, 0, 0, 0, 0, 0, 0, 0, 0),
                (29, 288, 32, 32, 69, 86, 192, 0, 0, 0, 0, 0, 0, 0, 0),
                (-180, 136, 154, 76, 32, 160, 32, 0, 0, 0, 0, 0, 0, 0, 0),
                (72, 32, 32, 32, 66, 32, 32, 0, 0, 0, 0, 0, 0, 0, 0),
                (887, 433, 38, 433, 64, 0, 205, 0, 0, 0, 0, 0, 0, -128, -128),
                (35, 242, 32, 288, 103, 73, 192, 0, 0, 0, 0, 0, 0, 0, 0),
                (131, -6, 32, 30, 248, 288, 245, 0, 0, 0, 0, 0, 0, 0, 0)
                );
    constant children_left : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 13, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 9, 3, 5, 7, -1, -1, -1, -1, 11, 13, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 13, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1)
                );
    constant children_right : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 14, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 10, 4, 6, 8, -1, -1, -1, -1, 12, 14, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 14, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1)
                );
    constant value_int : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((0, 0, 0, 0, 0, 0, 0, 3, -19, -20, -26, 26, 17, 4, -19),
                (0, 0, 0, 0, 0, 0, 0, 13, -9, -15, -21, 20, -11, 3, -15),
                (0, 0, 0, 0, 0, 0, 0, 3, -13, -19, -12, 19, 13, 3, -15),
                (0, 0, 0, 0, 0, 0, 0, 7, 16, -6, 7, -11, -17, 12, -9),
                (0, 0, 0, 0, 0, 0, 0, -10, 6, -15, -4, 15, 7, 0, -12),
                (0, 0, 0, 0, 0, 0, 0, 13, -8, 2, -10, -9, -15, 12, -5),
                (0, 0, 0, 0, 0, 0, 0, 7, -12, 10, -9, 10, -6, 0, -9),
                (0, 0, 0, 0, 0, 0, 0, 12, -2, -3, 6, 4, -9, -15, -9),
                (0, 0, 0, 0, 0, 0, 0, 8, -7, -1, -9, 0, -10, -10, -15),
                (0, 0, 0, 0, 0, 0, 0, -9, 3, -14, -2, 12, 8, 2, -9),
                (0, 0, 0, 0, 0, 0, 0, 9, -7, -2, 6, -4, -10, -13, -7),
                (0, 0, 0, 0, 0, 0, 0, 5, -4, -12, 8, -11, -3, 4, -9),
                (0, 0, 0, 0, 0, 0, 0, 11, 6, -2, 4, -13, 4, 0, -8),
                (0, 0, 0, 0, 0, 0, 0, -6, 3, 16, 6, -12, -6, -1, -8),
                (0, 0, 0, 0, 0, 0, 0, 5, -5, -8, -3, -10, -2, 7, 0),
                (0, 0, 0, 0, 0, 0, 0, 1, 8, -6, 2, -13, -8, 10, -5),
                (0, 0, 0, 0, 0, 0, 0, -6, 6, 11, 6, 0, -10, -7, -12),
                (0, 0, 0, 0, 0, 0, 0, 5, 17, -1, 4, -4, 2, 9, -3),
                (0, 0, 0, 0, 0, 0, 0, 7, 1, -10, 0, -14, -5, -3, -7),
                (0, 0, 0, 0, 0, 0, 0, 1, 8, -8, -3, -10, -4, 6, -2),
                (0, 0, 0, 0, 0, 0, 0, 2, -2, -9, 5, -17, -2, -12, -7),
                (0, 0, 0, 0, 0, 0, 0, 5, 15, 1, 6, -8, 0, -12, 4),
                (0, 0, 0, 0, 0, 0, 0, 3, 8, -9, 5, -12, 0, -11, 3),
                (0, 0, 0, 0, 0, 0, 0, 8, 3, 3, -1, -9, -13, -1, -11),
                (0, 0, 0, 0, 0, 0, 0, 1, -4, -7, -2, -10, -1, 12, -4),
                (0, 0, 0, 0, 0, 0, 0, 5, -8, 3, -2, 11, -2, 7, -3),
                (0, 0, 0, 0, 0, 0, 0, 2, 11, 5, 0, -9, -2, 2, -3),
                (0, 0, 0, 0, 0, 0, 0, -3, 1, 11, 1, -13, -6, -1, -9),
                (0, 0, 0, 0, 0, 0, 0, -9, 5, -9, 1, -14, -4, -5, -1),
                (0, 0, 0, 0, 0, 0, 0, 0, 2, -7, -1, -6, -1, 6, -1),
                (0, 0, 0, 0, 0, 0, 0, 3, -7, 2, -1, 9, -1, 0, -11),
                (0, 0, 0, 0, 0, 0, 0, 4, 12, 4, 0, 2, 9, -2, 1),
                (0, 0, 0, 0, 0, 0, 0, 7, -11, -7, 3, -9, 1, 4, -2),
                (0, 0, 0, 0, 0, 0, 0, -1, 1, -10, -2, -12, -3, -13, -7),
                (0, 0, 0, 0, 0, 0, 0, 3, 8, -10, 15, -1, 1, -5, -10),
                (0, 0, 0, 0, 0, 0, 0, -12, 0, 7, 2, -1, -10, 5, -2),
                (0, 0, 0, 0, 0, 0, 0, 8, 3, 0, -5, -7, -12, 5, -6),
                (0, 0, 0, 0, 0, 0, 0, -1, 1, -9, 3, -6, 0, 9, -7),
                (0, 0, 0, 0, 0, 0, 0, 8, -9, 2, -2, 1, -9, 5, -1),
                (0, 0, 0, 0, 0, 0, 0, -11, 2, -7, 0, -5, 3, -7, 0),
                (0, 0, 0, 0, 0, 0, 0, -1, 1, -11, -5, 13, 44, -12, 0),
                (0, 0, 0, 0, 0, 0, 0, -8, 0, 4, 0, -1, -5, 1, -6),
                (0, 0, 0, 0, 0, 0, 0, 2, -17, 0, -3, 10, 22, -13, 0),
                (0, 0, 0, 0, 0, 0, 0, -8, 3, 11, 6, 2, -16, -1, 1),
                (0, 0, 0, 0, 0, 0, 0, 3, 0, 4, -1, 1, -11, -2, -8),
                (0, 0, 0, 0, 0, 0, 0, -1, 0, 8, 0, -12, -6, 4, -7),
                (0, 0, 0, 0, 0, 0, 0, -2, 9, 8, -2, -1, 1, 3, -5),
                (0, 0, 0, 0, 0, 0, 9, -19, -11, 0, -2, -2, -8, 9, 9),
                (0, 0, 0, 0, 0, 0, 0, 5, 1, 2, -4, -1, 2, -2, 0),
                (0, 0, 0, 0, 0, 0, 0, 0, -7, -2, -9, 9, -1, -4, 3),
                (0, 0, 0, 0, 0, 0, 0, 9, 0, -1, -7, -2, 4, -6, 0),
                (0, 0, 0, 0, 0, 0, 0, 5, -6, 1, -3, 9, -4, -6, 1),
                (0, 0, 0, 0, 0, 0, 0, -2, 10, 12, 3, 0, 8, 0, -2),
                (0, 0, 0, 0, 0, 0, 0, -11, -1, -5, 1, -1, 3, -7, 0),
                (0, 0, 0, 0, 0, 0, 0, 7, 0, -3, 4, 3, 0, -6, 0),
                (0, 0, 0, 0, 0, 0, 0, -18, 12, -9, -17, 1, 0, -11, -3),
                (0, 0, 0, 0, 0, 0, 0, -1, 1, -1, -4, 3, -5, -3, -12),
                (0, 0, 0, 0, 0, 0, 0, -14, 14, -6, -16, 0, -7, -6, 1),
                (0, 0, 0, 0, 0, 0, 0, 13, 2, -1, -10, -1, 6, 0, -2),
                (0, 0, 0, 0, 0, 0, 0, -10, -3, 2, -3, 0, 1, -1, 1),
                (0, 0, 0, 0, 0, 0, 0, -7, 22, -4, 1, -3, 4, -7, 0),
                (0, 0, 0, 0, 0, 0, 0, -9, 1, 7, 0, 2, -1, -1, 5),
                (0, 0, 0, 0, 0, 0, 0, -8, 7, -8, -15, -3, 0, 4, 0),
                (0, 0, 0, 0, 0, 0, 0, 7, -12, 1, 6, -2, 0, 3, 0),
                (0, 0, 0, 0, 0, -13, 0, 0, 1, -2, 1, -4, -13, -13, -13),
                (0, 0, 0, 0, 0, 0, 0, -4, 7, 26, 6, 3, 0, -8, -1),
                (0, 0, 0, 0, 0, 0, 0, 6, -1, -23, 0, -11, 0, 2, -11),
                (0, 0, 0, 0, 0, 0, 0, -9, -1, 1, 7, -1, 2, 3, -3),
                (0, 0, 0, 0, 0, 0, 0, -5, 1, -3, 0, 5, -6, -4, 2),
                (0, 0, 0, 0, 0, 0, 0, 8, 13, -1, 2, 1, -1, -7, 0),
                (0, 0, 0, 0, 0, 0, 0, -14, -3, 0, -1, 4, 17, 6, -8),
                (0, 0, 0, 0, 0, 0, 0, -7, 7, 1, -1, -3, -11, 1, -6),
                (0, 0, 0, 0, 0, 0, 0, 1, -4, 3, 15, 0, 1, -5, 9),
                (0, 0, 0, 0, 0, 0, 0, 6, 0, -1, -9, -1, 3, -4, 0),
                (0, 0, 0, 0, 0, 0, 0, 3, -12, 3, 0, -4, 12, -14, -6),
                (0, 0, 0, 0, 0, 0, 0, 0, -8, 3, 0, 1, -8, 10, -2),
                (0, 0, 0, 0, 0, 0, 0, -6, 0, 2, -4, -4, -9, 2, -3),
                (0, 0, 0, 0, 0, 0, 0, 0, 5, -7, 1, 5, -5, -1, 2),
                (0, 0, 0, 0, 0, 0, 0, 0, -1, -11, -5, 5, -3, 14, 3),
                (0, 0, 0, 0, 0, 0, 0, 1, -4, -1, 7, 10, -7, -1, 0),
                (0, 0, 0, 0, 0, 0, 0, 2, -3, 1, 4, 1, 0, 0, -3),
                (0, 0, 0, 0, 0, 0, 0, 0, 4, -6, 0, -10, -1, 3, 0),
                (0, 0, 0, 0, 0, 0, 0, 3, 0, -2, -11, 8, 35, -2, 1),
                (0, 0, 0, 0, 0, 0, 0, -1, 1, 1, -2, -3, 2, 2, 6),
                (0, -14, 0, 0, 0, 1, 0, -1, 0, -14, -14, -14, -14, -14, -14),
                (0, 0, 0, 0, 0, 0, 0, 1, 0, -4, 3, -3, 10, -10, -3),
                (0, 0, 0, 0, 0, 0, 0, 6, -1, -2, 1, 2, 10, -15, 1),
                (0, 0, 0, 0, 0, 0, 0, -3, 1, 10, 2, 1, -4, -1, 0),
                (0, 0, 0, 0, 0, 0, 0, 15, -6, 0, 3, -2, 1, -10, -2),
                (0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 3, 7, -7, -5, 2),
                (0, 0, 0, 0, 0, 0, 0, 6, 0, 9, -2, 0, -2, 3, -3),
                (0, 0, 0, 0, 0, 0, 0, -2, 2, 0, -1, -10, 2, -4, -10),
                (0, 0, 0, 0, 0, 0, 0, 0, 5, 17, 3, 1, 9, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, 0, 5, 0, -1, -2, -9, 0, 7),
                (0, 0, 0, 0, 0, 0, 0, 0, -6, 3, -1, 0, 8, -1, 0),
                (0, 0, 0, 0, 0, 0, 0, 8, -6, 14, 8, -2, 0, -2, 1),
                (0, 0, 0, 0, 0, 0, 0, -6, 4, 5, 1, 0, 5, 0, -1),
                (0, 0, 0, 0, 0, 9, 0, 0, 13, -1, -11, -7, 3, 9, 9),
                (0, 0, 0, 0, 0, 0, 0, -2, 1, -1, -8, 0, 4, -1, 0),
                (0, 0, 0, 0, 0, 0, 0, 0, 2, 0, -1, -7, 3, -8, 10)
                );
    constant parent : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 6, 6, 5, 5),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 2, 2, 3, 3, 4, 4, 1, 1, 9, 9, 10, 10),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 6, 6, 5, 5),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6)
                );
    constant depth : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 3, 3, 3, 3, 2, 2, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3)
                );
    constant iLeaf : intArray2D(nTrees-1 downto 0)(nLeaves-1 downto 0) := ((7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (5, 6, 7, 8, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14)
                );
    constant value : tyArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := to_tyArray2D(value_int);
      constant threshold : txArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := to_txArray2D(threshold_int);
end Arrays0;