library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_misc.all;
  use ieee.numeric_std.all;

  use work.Constants.all;
  use work.Types.all;
  package Arrays0 is

    constant initPredict : ty := to_ty(0);
    constant feature : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((4, 1, 0, 3, 1, 0, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 1, 0, 0, 17, 3, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 4, 0, 3, 3, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 19, 0, 0, 15, 2, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 1, 3, 0, 3, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 3, 4, 17, 4, 18, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 16, 18, 18, 1, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 17, 5, 16, 4, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 16, 3, 4, 17, 16, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 7, 1, 17, 6, 5, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 0, 4, 3, 2, 5, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (7, 17, 6, 5, 12, 17, 13, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 3, 17, 20, 20, 7, 13, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 17, 1, 7, 14, 0, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 2, 1, 1, 16, 16, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 1, 16, 18, 16, 16, 10, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 10, 4, 1, 4, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 6, 14, 4, 7, 16, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 20, 17, 16, 16, 20, 12, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 1, 17, 3, 16, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 18, 4, 5, 4, 1, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 5, 19, 9, 4, 10, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 2, 1, 4, 3, 5, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 4, 4, 16, 16, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 16, 16, 0, 2, 17, 10, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 17, 3, 17, 13, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 7, 18, 13, 13, 16, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 4, 17, 16, 16, 5, 14, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 4, 4, 8, 2, 18, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 8, 2, 10, 5, 17, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 3, 12, 18, 17, 17, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 7, 14, 10, 11, 15, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 4, 10, 0, 2, 20, 8, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 17, 1, 5, 9, 4, 19, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 18, 16, 19, 4, 19, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 16, 17, 0, 2, 16, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 20, 15, 13, 16, 12, 13, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 2, 17, 4, 16, 5, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 2, 18, 4, 3, 3, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 6, 6, 16, 17, 20, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 17, 0, 16, 16, 17, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 2, 16, -2, 16, 2, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 16, 17, 2, 10, 18, 19, -2, -2, -2, -2, -2, -2, -2, -2),
                (19, 11, 17, 17, 2, 4, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 16, 4, 1, 1, 1, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 3, 19, 9, 4, 16, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (19, 9, 17, 10, 16, 20, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 4, 0, 1, 16, 1, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 13, 1, 5, 3, 4, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 6, 2, 18, 0, 1, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (8, 10, 5, 17, 5, 9, 9, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 18, 6, 17, 17, 0, 20, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 10, 1, 17, 0, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 16, 16, 4, 16, 2, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 17, 17, 4, 2, 2, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 1, 15, 1, 3, 16, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 17, -2, 17, 16, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 16, 10, 4, 4, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 17, 0, 4, 12, -2, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 18, 6, 3, 18, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 5, 4, 2, 2, 16, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 3, 19, 17, 17, 3, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 4, 19, 16, 16, 20, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 0, 8, 3, 9, 20, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 1, 17, 2, -2, 17, 19, -2, -2, -2, -2, -2, -2, -2, -2),
                (11, 17, 7, 17, 17, 14, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 9, 4, 20, 16, 8, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 17, 2, 17, 15, 2, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 3, 3, 9, 17, 4, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 4, 0, 11, 16, 17, 15, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 17, 2, 3, 2, 16, 14, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 7, 0, 17, 5, 2, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 20, 11, 6, 3, 17, 19, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 0, 2, 17, 12, 4, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 1, 10, 2, 4, 17, 9, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 5, 16, 16, 16, 16, 5, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 4, 0, 17, 18, 17, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 5, 17, 2, 7, 0, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 0, 12, 16, 0, 3, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 1, 1, 1, 4, 1, 19, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 18, 3, 17, 17, 1, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 17, 4, 3, 13, 18, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 3, 2, 2, 17, -2, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 1, 16, 0, 18, 3, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 20, 20, 20, 0, 10, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (20, 12, 17, 3, 4, 17, 12, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 16, 17, 0, 2, 13, 15, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 9, 4, 19, 8, 2, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 3, 1, 3, 0, 17, 6, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 20, 0, 16, 20, 14, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 3, 1, 18, 18, 1, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 15, 3, 17, 17, 17, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 0, 16, 0, 1, 1, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 16, 0, 2, 1, 20, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 15, 14, 20, 17, 15, 3, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 6, 16, 11, 17, 17, 20, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 4, 2, 9, 1, 0, 7, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 4, 16, 17, 0, 18, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 1, 1, 1, 16, 3, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 17, 2, 17, 16, 1, 3, -2, -2, -2, -2, -2, -2, -2, -2)
                );
    constant threshold_int : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((288, 29, 215, 89, 59, 175, 130, 0, 0, 0, 0, 0, 0, 0, 0),
                (288, 18, 238, 163, 205, 143, 35, 0, 0, 0, 0, 0, 0, 0, 0),
                (49, 189, 352, 136, 121, 89, 286, 0, 0, 0, 0, 0, 0, 0, 0),
                (288, 160, 170, 104, 32, 72, 352, 0, 0, 0, 0, 0, 0, 0, 0),
                (70, 291, 91, 134, 363, 91, 160014, 0, 0, 0, 0, 0, 0, 0, 0),
                (542, 112, 352, 200, 352, 696, 154, 0, 0, 0, 0, 0, 0, 0, 0),
                (80, 151, 134904, 711, 471, 108, 67, 0, 0, 0, 0, 0, 0, 0, 0),
                (6, 317, 53, 32, 11658, 352, 79, 0, 0, 0, 0, 0, 0, 0, 0),
                (352, 79266, 154, 288, 199, 87466, 240, 0, 0, 0, 0, 0, 0, 0, 0),
                (127, 32, 100, 142, 32, 32, 124, 0, 0, 0, 0, 0, 0, 0, 0),
                (628, 387, 288, 162, 427, 32, 150, 0, 0, 0, 0, 0, 0, 0, 0),
                (32, 146, 32, 32, 32, 65, 32, 0, 0, 0, 0, 0, 0, 0, 0),
                (36, 128, 231, 288, 288, 32, 32, 0, 0, 0, 0, 0, 0, 0, 0),
                (100, 128, 106, 32, 32, 284, 171227, 0, 0, 0, 0, 0, 0, 0, 0),
                (85, -32, -18, 126, 25440, 139086, 347, 0, 0, 0, 0, 0, 0, 0, 0),
                (343, 119, 6883, 816, 158482, 6175, 32, 0, 0, 0, 0, 0, 0, 0, 0),
                (38, 32, 352, 32, 288, 65040, 70243, 0, 0, 0, 0, 0, 0, 0, 0),
                (277, 32, 32, 288, 32, 46598, 148, 0, 0, 0, 0, 0, 0, 0, 0),
                (26, 288, 137, 186326, 144767, 160, 32, 0, 0, 0, 0, 0, 0, 0, 0),
                (412, 127, 96, 181, 183165, 18343, 16219, 0, 0, 0, 0, 0, 0, 0, 0),
                (186886, 771, 288, 32, 288, 15, 276, 0, 0, 0, 0, 0, 0, 0, 0),
                (46, 32, 96, 32, 352, 32, 138, 0, 0, 0, 0, 0, 0, 0, 0),
                (1861, 163, -56, 288, 112, 32, -33, 0, 0, 0, 0, 0, 0, 0, 0),
                (287, 288, 288, 91121, 124283, 119837, 127708, 0, 0, 0, 0, 0, 0, 0, 0),
                (381, 14226, 10077, 226, 233, 95, 32, 0, 0, 0, 0, 0, 0, 0, 0),
                (-33, 101, 228, 62, 32, 1498, 144618, 0, 0, 0, 0, 0, 0, 0, 0),
                (135, 32, 178, 32, 32, 109234, 402, 0, 0, 0, 0, 0, 0, 0, 0),
                (70, 288, 121, 147813, 39584, 32, 32, 0, 0, 0, 0, 0, 0, 0, 0),
                (155881, 352, 288, 32, 180, 414, 130, 0, 0, 0, 0, 0, 0, 0, 0),
                (37, 32, 208, 32, 32, 93, 34018, 0, 0, 0, 0, 0, 0, 0, 0),
                (49, -308, 32, 139, 94, 172, 192, 0, 0, 0, 0, 0, 0, 0, 0),
                (166, 32, 32, 32, 32, 32, 288, 0, 0, 0, 0, 0, 0, 0, 0),
                (16499, 288, 32, 115, 286, 288, 32, 0, 0, 0, 0, 0, 0, 0, 0),
                (186359, 93, 36, 32, 32, 288, 96, 0, 0, 0, 0, 0, 0, 0, 0),
                (149, 902, 119788, 96, 352, 288, 189, 0, 0, 0, 0, 0, 0, 0, 0),
                (139, 2618, 144, 204, 427, 184663, 39, 0, 0, 0, 0, 0, 0, 0, 0),
                (149, 160, 32, 32, 99502, 32, 32, 0, 0, 0, 0, 0, 0, 0, 0),
                (66, 249, 85, 288, 97461, 32, 72, 0, 0, 0, 0, 0, 0, 0, 0),
                (100, 70, 358, 288, 120, 5, 542, 0, 0, 0, 0, 0, 0, 0, 0),
                (228, 32, 32, 100540, 188, 288, -92, 0, 0, 0, 0, 0, 0, 0, 0),
                (-100, 92, -6, 131281, 44507, 9, 369, 0, 0, 0, 0, 0, 0, 0, 0),
                (-134, -347, 18277, 0, 101379, 166, 239, 0, 0, 0, 0, 0, 0, -128, -128),
                (242, 3655, 279, 202, 32, 456, 288, 0, 0, 0, 0, 0, 0, 0, 0),
                (96, 32, 120, 101, 307, 352, -22, 0, 0, 0, 0, 0, 0, 0, 0),
                (183033, 159948, 288, 106, 50, 15, 150, 0, 0, 0, 0, 0, 0, 0, 0),
                (148, 130, 288, 32, 288, 93805, -4, 0, 0, 0, 0, 0, 0, 0, 0),
                (96, 32, 125, 32, 65468, 96, 157, 0, 0, 0, 0, 0, 0, 0, 0),
                (78, 288, 99, 18, 56247, -48, 340, 0, 0, 0, 0, 0, 0, 0, 0),
                (-43, 32, 17, 32, 106, 288, 75643, 0, 0, 0, 0, 0, 0, 0, 0),
                (-30, 32, 434, 81, -153, 139, 21, 0, 0, 0, 0, 0, 0, 0, 0),
                (32, 32, 32, 101, 32, 32, 32, 0, 0, 0, 0, 0, 0, 0, 0),
                (729, 546, 32, 238, 195, 187, 96, 0, 0, 0, 0, 0, 0, 0, 0),
                (-13, 32, -11, 65, 284, 183626, 100474, 0, 0, 0, 0, 0, 0, 0, 0),
                (239, 26543, 5302, 288, 134410, 239, 147138, 0, 0, 0, 0, 0, 0, 0, 0),
                (187330, 5, 132, 288, -33, 44, 142, 0, 0, 0, 0, 0, 0, 0, 0),
                (64, 50, 32, 41, 93, 101346, 272, 0, 0, 0, 0, 0, 0, 0, 0),
                (-267, 142, 100, 0, 100, 107933, 171, 0, 0, 0, 0, 0, 0, -128, -128),
                (259, 31911, 32, 288, 288, 46532, 96868, 0, 0, 0, 0, 0, 0, 0, 0),
                (59, 64, 59, 288, 32, 0, 1, 0, 0, 0, 0, 0, 0, -128, -128),
                (913, 13, 32, 150, 21, 136517, 26576, 0, 0, 0, 0, 0, 0, 0, 0),
                (223, 32, 288, 99, 99, 59672, 456, 0, 0, 0, 0, 0, 0, 0, 0),
                (669, 226, 160, 101, 282, 205, -79, 0, 0, 0, 0, 0, 0, 0, 0),
                (239, 288, 288, 106204, 56049, 32, 147, 0, 0, 0, 0, 0, 0, 0, 0),
                (120, 197, 32, 79, 32, 160, 187, 0, 0, 0, 0, 0, 0, 0, 0),
                (971, 30, 234, 302, 0, 233, 160, 0, 0, 0, 0, 0, 0, -128, -128),
                (32, 102, 32, 69, 165, 32, 288, 0, 0, 0, 0, 0, 0, 0, 0),
                (77, 32, 352, 288, 80204, 32, 181, 0, 0, 0, 0, 0, 0, 0, 0),
                (271, 254, 200, 254, 32, 86, 37361, 0, 0, 0, 0, 0, 0, 0, 0),
                (-44, -240, 13, 32, 8, 288, 19, 0, 0, 0, 0, 0, 0, 0, 0),
                (157, 352, 180, 32, 56280, 153, 32, 0, 0, 0, 0, 0, 0, 0, 0),
                (321, 312, 341, 120, 321, 125123, 32, 0, 0, 0, 0, 0, 0, 0, 0),
                (90, 32, 96, 197, 32, 70, 45989, 0, 0, 0, 0, 0, 0, 0, 0),
                (136, 160, 32, 32, 164, 164, 160, 0, 0, 0, 0, 0, 0, 0, 0),
                (180464, 239, 217, 94, 32, 288, 57, 0, 0, 0, 0, 0, 0, 0, 0),
                (17, 0, 32, 319, 288, 106, 32, 0, 0, 0, 0, 0, 0, 0, 0),
                (263, 32, 156276, 65023, 59178, 6175, 32, 0, 0, 0, 0, 0, 0, 0, 0),
                (114, 288, 123, 322, 92, 6, 124, 0, 0, 0, 0, 0, 0, 0, 0),
                (73, 32, 84, 130, 32, 382, 128894, 0, 0, 0, 0, 0, 0, 0, 0),
                (144, 154, 32, 10769, 154, -39, 155, 0, 0, 0, 0, 0, 0, 0, 0),
                (239, 39, 35, 18, 288, 23, 288, 0, 0, 0, 0, 0, 0, 0, 0),
                (-308, 246, -217, 83, 123, 33, -179, 0, 0, 0, 0, 0, 0, 0, 0),
                (291, 203, 288, 193, 32, 411, 437, 0, 0, 0, 0, 0, 0, 0, 0),
                (3622, 57, -394, 144, 197, 0, -180, 0, 0, 0, 0, 0, 0, -128, -128),
                (366, 91, 130639, 93, 84, -9, 102, 0, 0, 0, 0, 0, 0, 0, 0),
                (59836, 352, 352, 32, 318, 32, 53, 0, 0, 0, 0, 0, 0, 0, 0),
                (32, 32, 273, 190, 288, 270, 32, 0, 0, 0, 0, 0, 0, 0, 0),
                (239, 6734, 190, 197, 234, 32, 32, 0, 0, 0, 0, 0, 0, 0, 0),
                (71, 32, 352, 96, 32, 307, 313, 0, 0, 0, 0, 0, 0, 0, 0),
                (130, 128, 49, 128, 265, 237, 32, 0, 0, 0, 0, 0, 0, 0, 0),
                (123, 96, 132, 187594, 160, 32, -22, 0, 0, 0, 0, 0, 0, 0, 0),
                (9, 80, 29, 422, 36, 28, 129223, 0, 0, 0, 0, 0, 0, 0, 0),
                (-52, 32, -52, 126, 256, 88, -52, 0, 0, 0, 0, 0, 0, 0, 0),
                (362, 358, 115984, 356, -2, 72, 151, 0, 0, 0, 0, 0, 0, 0, 0),
                (146611, 145409, 338, 288, 25, 288, 388, 0, 0, 0, 0, 0, 0, 0, 0),
                (203, 32, 32, 96, 176, 32, 32, 0, 0, 0, 0, 0, 0, 0, 0),
                (71, 32, 98580, 32, 249, 8, 352, 0, 0, 0, 0, 0, 0, 0, 0),
                (154, 288, 84, 32, 85, 219, 32, 0, 0, 0, 0, 0, 0, 0, 0),
                (5170, 288, 6685, 75, 208, 163, 440, 0, 0, 0, 0, 0, 0, 0, 0),
                (49, 48, 56, 48, 125814, 123, 4, 0, 0, 0, 0, 0, 0, 0, 0),
                (25, 322, 25, 204, 187232, -16, 120, 0, 0, 0, 0, 0, 0, 0, 0)
                );
    constant children_left : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 13, 7, 9, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 13, 7, 9, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 13, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 13, 9, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 13, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1)
                );
    constant children_right : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 14, 8, 10, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 14, 8, 10, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 14, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 14, 10, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 14, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1)
                );
    constant value_int : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((0, 0, 0, 0, 0, 0, 0, 7, -37, -38, -54, 53, 34, 9, -40),
                (0, 0, 0, 0, 0, 0, 0, 30, -14, -35, -14, 33, -18, 3, -27),
                (0, 0, 0, 0, 0, 0, 0, 31, 19, 4, -22, -21, -33, 19, -12),
                (0, 0, 0, 0, 0, 0, 0, 14, -22, 23, -14, 28, 21, -8, 11),
                (0, 0, 0, 0, 0, 0, 0, 15, -14, -5, -21, -8, -23, -29, -16),
                (0, 0, 0, 0, 0, 0, 0, 4, 21, -18, 3, -21, -31, 12, -26),
                (0, 0, 0, 0, 0, 0, 0, 16, -20, 1, -14, -19, -28, 0, -16),
                (0, 0, 0, 0, 0, 0, 0, 19, 6, -28, -3, -21, 8, 4, -9),
                (0, 0, 0, 0, 0, 0, 0, -20, 1, -3, 13, 16, 3, -6, -22),
                (0, 0, 0, 0, 0, 0, 0, -27, 9, -17, 19, 8, -3, -16, -25),
                (0, 0, 0, 0, 0, 0, 0, 3, -12, -14, -26, -15, -25, 15, -6),
                (0, 0, 0, 0, 0, 0, 0, 6, -31, -22, 7, -21, -4, 8, -6),
                (0, 0, 0, 0, 0, 0, 0, 11, 19, -13, 14, -9, 0, -20, 8),
                (0, 0, 0, 0, 0, 0, 0, -19, 2, 11, 1, -1, -8, -22, 1),
                (0, 0, 0, 0, 0, 0, 0, 19, -17, 26, 6, 5, -1, 0, -7),
                (0, 0, 0, 0, 0, 0, 0, 1, -16, -20, -1, -33, -20, -3, -14),
                (0, 0, 0, 0, 0, 0, 0, 2, 10, -22, 0, -8, -1, 10, -3),
                (0, 0, 0, 0, 0, 0, 0, -12, 1, -3, 2, -23, 21, 4, -8),
                (0, 0, 0, 0, 0, 0, 0, 2, 31, 20, 7, -15, -1, -12, 4),
                (0, 0, 0, 0, 0, 0, 0, 1, -7, -18, 17, -6, -26, -30, -7),
                (0, 0, 0, 0, 0, 0, 0, 3, -1, -15, -1, 19, 46, -3, -33),
                (0, 0, 0, 0, 0, 0, 0, -19, 17, -10, 1, 9, -4, -6, 1),
                (0, 0, 0, 0, 0, 0, 0, -27, 21, -39, -18, 11, 2, 4, -1),
                (0, 0, 0, 0, 0, 0, 0, -6, 10, 3, -7, -10, 0, 5, -5),
                (0, 0, 0, 0, 0, 0, 0, 21, -12, -1, 2, -10, -28, -2, -10),
                (0, 0, 0, 0, 0, 0, 0, 7, 21, -16, 6, -30, 0, -14, 4),
                (0, 0, 0, 0, 0, 0, 0, -10, 2, 2, -5, -18, 2, -21, 28),
                (0, 0, 0, 0, 0, 0, 0, -11, 3, 24, 7, 5, -3, 4, -2),
                (0, 0, 0, 0, 0, 0, 0, -2, 2, 8, 0, 7, -4, -8, 5),
                (0, 0, 0, 0, 0, 0, 0, -1, -19, 8, -3, 5, -4, -5, 2),
                (0, 0, 0, 0, 0, 0, 0, -101, 2, 13, 4, 0, -15, -3, 2),
                (0, 0, 0, 0, 0, 0, 0, -9, 6, -1, 3, 20, -12, -5, 2),
                (0, 0, 0, 0, 0, 0, 0, 14, -15, 19, -4, 1, -6, -18, -1),
                (0, 0, 0, 0, 0, 0, 0, 8, 0, 0, -8, 10, -1, 34, 10),
                (0, 0, 0, 0, 0, 0, 0, 1, -1, -17, 17, -6, -17, -11, 3),
                (0, 0, 0, 0, 0, 0, 0, 4, -26, 0, -8, -23, 0, 7, -14),
                (0, 0, 0, 0, 0, 0, 0, 3, -14, 2, -1, -8, 5, -13, 1),
                (0, 0, 0, 0, 0, 0, 0, -4, 3, 0, -22, 18, 5, 1, -2),
                (0, 0, 0, 0, 0, 0, 0, -3, 6, 0, 2, 12, -4, -15, -6),
                (0, 0, 0, 0, 0, 0, 0, -6, 1, 0, 3, -3, 67, 9, -17),
                (0, 0, 0, 0, 0, 0, 0, 14, 2, -13, 3, -24, 16, 0, 36),
                (0, 0, 0, -54, 0, 0, 0, -4, 16, 16, -2, -1, 1, -54, -54),
                (0, 0, 0, 0, 0, 0, 0, 7, -25, 0, -1, -16, 0, 12, -10),
                (0, 0, 0, 0, 0, 0, 0, 0, -5, 6, 23, -9, 3, 4, 0),
                (0, 0, 0, 0, 0, 0, 0, 0, -5, -3, 5, 4, 16, -4, 15),
                (0, 0, 0, 0, 0, 0, 0, 1, -1, -4, 8, -5, 2, -20, -1),
                (0, 0, 0, 0, 0, 0, 0, 8, -11, 3, -2, 55, -3, -2, 1),
                (0, 0, 0, 0, 0, 0, 0, -8, 1, 16, 5, -39, -10, 0, -2),
                (0, 0, 0, 0, 0, 0, 0, 12, 1, 0, -4, -4, 0, -3, 2),
                (0, 0, 0, 0, 0, 0, 0, 24, -18, -24, 27, 0, -11, 15, -10),
                (0, 0, 0, 0, 0, 0, 0, 8, 0, -24, -4, -17, 8, 5, -1),
                (0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 8, -2, 14, 9, -8),
                (0, 0, 0, 0, 0, 0, 0, -7, 1, 5, -3, -4, -25, -1, 0),
                (0, 0, 0, 0, 0, 0, 0, -11, 13, -3, 0, 26, -18, 1, -2),
                (0, 0, 0, 0, 0, 0, 0, -10, 1, 3, 0, 34, 9, -28, 1),
                (0, 0, 0, 0, 0, 0, 0, 0, -3, 6, -2, -3, 2, -13, 2),
                (0, 0, 0, 0, 0, 0, 0, 0, -54, 2, -1, -2, 0, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, -10, 11, 2, -1, -3, 1, -2, -12),
                (0, 0, 0, 0, 0, -63, 0, -9, 11, 12, -1, 7, 0, -63, -63),
                (0, 0, 0, 0, 0, 0, 0, -1, -10, 3, 0, -5, 31, 25, -14),
                (0, 0, 0, 0, 0, 0, 0, -7, 4, 3, 0, -7, -1, -1, 5),
                (0, 0, 0, 0, 0, 0, 0, 1, 0, -8, 4, -6, 18, -18, 4),
                (0, 0, 0, 0, 0, 0, 0, -5, 4, 6, -3, -7, 0, 7, -8),
                (0, 0, 0, 0, 0, 0, 0, -1, 3, 0, -3, 1, -8, 0, 7),
                (0, 0, 0, 0, 0, 0, 0, -38, -5, 0, 17, 13, -1, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, 0, 2, -10, 0, -4, 1, 5, 1),
                (0, 0, 0, 0, 0, 0, 0, 1, 12, 2, -3, -3, 1, 6, -1),
                (0, 0, 0, 0, 0, 0, 0, 0, 16, 4, -9, 5, -5, -10, 4),
                (0, 0, 0, 0, 0, 0, 0, 4, -35, -9, 25, 1, -4, 4, 0),
                (0, 0, 0, 0, 0, 0, 0, -1, -8, 12, 1, 2, 8, 0, -1),
                (0, 0, 0, 0, 0, 0, 0, 0, 1, -2, -15, 10, 0, 7, -15),
                (0, 0, 0, 0, 0, 0, 0, 11, -3, -13, 1, -2, -16, -1, 0),
                (0, 0, 0, 0, 0, 0, 0, 23, -6, 0, -4, -10, 0, 9, 0),
                (0, 0, 0, 0, 0, 0, 0, 0, -2, -1, 2, 7, 1, -25, -1),
                (0, 0, 0, 0, 0, 0, 0, 0, 3, -5, 0, 3, 0, -10, 0),
                (0, 0, 0, 0, 0, 0, 0, -12, 5, 3, -1, -12, 0, -11, -2),
                (0, 0, 0, 0, 0, 0, 0, -3, 17, -1, 6, -27, -4, 12, 0),
                (0, 0, 0, 0, 0, 0, 0, -7, 11, -8, -1, 5, -11, -1, 1),
                (0, 0, 0, 0, 0, 0, 0, 17, 0, -49, 0, 0, -18, -10, 10),
                (0, 0, 0, 0, 0, 0, 0, 0, 3, 0, -6, 0, -3, 1, 10),
                (0, 0, 0, 0, 0, 0, 0, 12, -39, -6, 35, 5, 21, -9, 0),
                (0, 0, 0, 0, 0, 0, 0, 1, -7, -8, 0, 0, -3, -1, 2),
                (0, 0, 0, 0, 0, -40, 0, 0, -26, -5, 26, 8, 0, -40, -40),
                (0, 0, 0, 0, 0, 0, 0, 2, 0, 4, -3, -29, 9, 40, 0),
                (0, 0, 0, 0, 0, 0, 0, 9, -2, 8, -1, 0, 3, -7, -1),
                (0, 0, 0, 0, 0, 0, 0, 20, 125, -7, 2, 0, -8, -16, 3),
                (0, 0, 0, 0, 0, 0, 0, 15, -7, 0, -9, 1, -3, 6, -1),
                (0, 0, 0, 0, 0, 0, 0, 4, 0, 4, -1, -2, 1, 2, -3),
                (0, 0, 0, 0, 0, 0, 0, 0, 13, -9, -1, 4, -2, 2, -5),
                (0, 0, 0, 0, 0, 0, 0, 48, -23, -6, 0, -8, 0, 4, 0),
                (0, 0, 0, 0, 0, 0, 0, -3, -13, -10, 2, 0, -7, -1, 2),
                (0, 0, 0, 0, 0, 0, 0, -3, 4, -18, 3, -3, 34, -57, 0),
                (0, 0, 0, 0, 0, 0, 0, 0, 7, 2, -9, 3, -5, -10, 16),
                (0, 0, 0, 0, 0, 0, 0, 0, 1, 10, 0, 0, -3, -10, 8),
                (0, 0, 0, 0, 0, 0, 0, 6, 0, 12, 1, 9, -7, -6, -1),
                (0, 0, 0, 0, 0, 0, 0, -6, 0, 1, -13, 3, -2, 1, -2),
                (0, 0, 0, 0, 0, 0, 0, -4, 2, 2, 17, -10, 5, -1, 0),
                (0, 0, 0, 0, 0, 0, 0, -26, 0, 19, -9, -1, 14, 0, -7),
                (0, 0, 0, 0, 0, 0, 0, 0, 11, -11, -1, 5, -4, -6, 0),
                (0, 0, 0, 0, 0, 0, 0, 2, -5, 19, -60, -45, 2, 0, 0)
                );
    constant parent : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 4, 4, 5, 5, 6, 6, 3, 3),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 4, 4, 5, 5, 6, 6, 3, 3),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 6, 6, 5, 5),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 5, 5, 6, 6, 4, 4),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 6, 6, 5, 5),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6)
                );
    constant depth : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3)
                );
    constant iLeaf : intArray2D(nTrees-1 downto 0)(nLeaves-1 downto 0) := ((7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14)
                );
    constant value : tyArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := to_tyArray2D(value_int);
      constant threshold : txArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := to_txArray2D(threshold_int);
end Arrays0;